
/////////////////////////////////////////////////////////////////
// Constants Define
/////////////////////////////////////////////////////////////////

`define MAP_WALL    3'b010
`define MAP_ROAD0   3'b000
`define MAP_ROAD1   3'b001
`define MAP_STAIRS  3'b011

/////////////////////////////////////////////////////////////////
// Constants Define
/////////////////////////////////////////////////////////////////

module mt(input clk,
		  input rst,
		  input sw_map,
		  input [5:0] gen_map_x1,
		  input [5:0] gen_map_y1,
		  output [2:0] gen_map_return1,
		  
		  input [5:0] gen_map_x2,
		  input [5:0] gen_map_y2,
		  output [2:0] gen_map_return2
);

	reg [2:0] mt [0:9] [0:19];
	
	assign gen_map_return1 = mt[gen_map_y1][gen_map_x1];
	assign gen_map_return2 = mt[gen_map_y2][gen_map_x2];
	
	parameter S0_RESET = 3'b000;
	parameter S1_MAP01 = 3'b001;
	/*parameter S2_SLI = 3'b010;
	parameter S3_BOX = 3'b011;
	parameter S4_SPL = 3'b100;*/
	reg [2:0] state, next_state;
	
	always @(posedge clk) begin
		if (rst == 1'b1) begin
			state = S0_RESET;
		end
		else begin
			state = next_state;
		end
		
		case (state)
			S0_RESET: begin
				
			end
			S1_MAP01: begin
				mt[0][0] = 3'b010;
				mt[0][1] = 3'b010;
				mt[0][2] = 3'b010;
				mt[0][3] = 3'b010;
				mt[0][4] = 3'b010;
				mt[0][5] = 3'b010;
				mt[0][6] = 3'b010;
				mt[0][7] = 3'b010;
				mt[0][8] = 3'b010;
				mt[0][9] = 3'b010;
				mt[0][10] = 3'b010;
				mt[0][11] = 3'b010;
				mt[0][12] = 3'b010;
				mt[0][13] = 3'b010;
				mt[0][14] = 3'b010;
				mt[0][15] = 3'b010;
				mt[0][16] = 3'b010;
				mt[0][17] = 3'b010;
				mt[0][18] = 3'b010;
				mt[0][19] = 3'b010;
				
				mt[1][0] = 3'b010;
				mt[1][1] = 3'b000;
				mt[1][2] = 3'b001;
				mt[1][3] = 3'b001;
				mt[1][4] = 3'b010;
				mt[1][5] = 3'b010;
				mt[1][6] = 3'b010;
				mt[1][7] = 3'b001;
				mt[1][8] = 3'b010;
				mt[1][9] = 3'b010;
				mt[1][10] = 3'b000;
				mt[1][11] = 3'b000;
				mt[1][12] = 3'b001;
				mt[1][13] = 3'b000;
				mt[1][14] = 3'b000;
				mt[1][15] = 3'b001;
				mt[1][16] = 3'b001;
				mt[1][17] = 3'b000;
				mt[1][18] = 3'b000;
				mt[1][19] = 3'b010;
				
				mt[2][0] = 3'b010;
				mt[2][1] = 3'b000;
				mt[2][2] = 3'b010;
				mt[2][3] = 3'b000;
				mt[2][4] = 3'b010;
				mt[2][5] = 3'b010;
				mt[2][6] = 3'b010;
				mt[2][7] = 3'b001;
				mt[2][8] = 3'b001;
				mt[2][9] = 3'b000;
				mt[2][10] = 3'b000;
				mt[2][11] = 3'b010;
				mt[2][12] = 3'b010;
				mt[2][13] = 3'b010;
				mt[2][14] = 3'b011;
				mt[2][15] = 3'b010;
				mt[2][16] = 3'b010;
				mt[2][17] = 3'b010;
				mt[2][18] = 3'b000;
				mt[2][19] = 3'b010;
				
				mt[3][0] = 3'b010;
				mt[3][1] = 3'b001;
				mt[3][2] = 3'b010;
				mt[3][3] = 3'b000;
				mt[3][4] = 3'b000;
				mt[3][5] = 3'b001;
				mt[3][6] = 3'b000;
				mt[3][7] = 3'b010;
				mt[3][8] = 3'b000;
				mt[3][9] = 3'b010;
				mt[3][10] = 3'b010;
				mt[3][11] = 3'b010;
				mt[3][12] = 3'b010;
				mt[3][13] = 3'b010;
				mt[3][14] = 3'b010;
				mt[3][15] = 3'b010;
				mt[3][16] = 3'b001;
				mt[3][17] = 3'b001;
				mt[3][18] = 3'b000;
				mt[3][19] = 3'b010;
				
				mt[4][0] = 3'b010;
				mt[4][1] = 3'b001;
				mt[4][2] = 3'b010;
				mt[4][3] = 3'b001;
				mt[4][4] = 3'b010;
				mt[4][5] = 3'b000;
				mt[4][6] = 3'b010;
				mt[4][7] = 3'b010;
				mt[4][8] = 3'b000;
				mt[4][9] = 3'b010;
				mt[4][10] = 3'b010;
				mt[4][11] = 3'b010;
				mt[4][12] = 3'b010;
				mt[4][13] = 3'b000;
				mt[4][14] = 3'b000;
				mt[4][15] = 3'b001;
				mt[4][16] = 3'b001;
				mt[4][17] = 3'b010;
				mt[4][18] = 3'b010;
				mt[4][19] = 3'b010;
				
				mt[5][0] = 3'b010;
				mt[5][1] = 3'b010;
				mt[5][2] = 3'b010;
				mt[5][3] = 3'b010;
				mt[5][4] = 3'b010;
				mt[5][5] = 3'b001;
				mt[5][6] = 3'b001;
				mt[5][7] = 3'b000;
				mt[5][8] = 3'b000;
				mt[5][9] = 3'b000;
				mt[5][10] = 3'b000;
				mt[5][11] = 3'b001;
				mt[5][12] = 3'b001;
				mt[5][13] = 3'b000;
				mt[5][14] = 3'b010;
				mt[5][15] = 3'b010;
				mt[5][16] = 3'b001;
				mt[5][17] = 3'b001;
				mt[5][18] = 3'b000;
				mt[5][19] = 3'b010;
				
				mt[6][0] = 3'b010;
				mt[6][1] = 3'b000;
				mt[6][2] = 3'b010;
				mt[6][3] = 3'b001;
				mt[6][4] = 3'b000;
				mt[6][5] = 3'b001;
				mt[6][6] = 3'b001;
				mt[6][7] = 3'b010;
				mt[6][8] = 3'b001;
				mt[6][9] = 3'b010;
				mt[6][10] = 3'b010;
				mt[6][11] = 3'b010;
				mt[6][12] = 3'b010;
				mt[6][13] = 3'b001;
				mt[6][14] = 3'b010;
				mt[6][15] = 3'b010;
				mt[6][16] = 3'b010;
				mt[6][17] = 3'b010;
				mt[6][18] = 3'b000;
				mt[6][19] = 3'b010;
				
				mt[7][0] = 3'b010;
				mt[7][1] = 3'b001;
				mt[7][2] = 3'b010;
				mt[7][3] = 3'b000;
				mt[7][4] = 3'b010;
				mt[7][5] = 3'b010;
				mt[7][6] = 3'b000;
				mt[7][7] = 3'b010;
				mt[7][8] = 3'b000;
				mt[7][9] = 3'b001;
				mt[7][10] = 3'b010;
				mt[7][11] = 3'b010;
				mt[7][12] = 3'b000;
				mt[7][13] = 3'b000;
				mt[7][14] = 3'b000;
				mt[7][15] = 3'b000;
				mt[7][16] = 3'b001;
				mt[7][17] = 3'b010;
				mt[7][18] = 3'b001;
				mt[7][19] = 3'b010;
				
				mt[8][0] = 3'b010;
				mt[8][1] = 3'b000;
				mt[8][2] = 3'b000;
				mt[8][3] = 3'b000;
				mt[8][4] = 3'b010;
				mt[8][5] = 3'b010;
				mt[8][6] = 3'b000;
				mt[8][7] = 3'b010;
				mt[8][8] = 3'b010;
				mt[8][9] = 3'b000;
				mt[8][10] = 3'b001;
				mt[8][11] = 3'b001;
				mt[8][12] = 3'b000;
				mt[8][13] = 3'b010;
				mt[8][14] = 3'b010;
				mt[8][15] = 3'b010;
				mt[8][16] = 3'b000;
				mt[8][17] = 3'b000;
				mt[8][18] = 3'b000;
				mt[8][19] = 3'b010;
				
				mt[9][0] = 3'b010;
				mt[9][1] = 3'b010;
				mt[9][2] = 3'b010;
				mt[9][3] = 3'b010;
				mt[9][4] = 3'b010;
				mt[9][5] = 3'b010;
				mt[9][6] = 3'b010;
				mt[9][7] = 3'b010;
				mt[9][8] = 3'b010;
				mt[9][9] = 3'b010;
				mt[9][10] = 3'b010;
				mt[9][11] = 3'b010;
				mt[9][12] = 3'b010;
				mt[9][13] = 3'b010;
				mt[9][14] = 3'b010;
				mt[9][15] = 3'b010;
				mt[9][16] = 3'b010;
				mt[9][17] = 3'b010;
				mt[9][18] = 3'b010;
				mt[9][19] = 3'b010;
				
			end
		endcase
	end
	
	always @* begin
		next_state = S0_RESET;
		case (state)
			S0_RESET: begin
				if (sw_map == 1) begin
					next_state = S1_MAP01;
				end /*else if (btnR == 1) begin
					next_state = S2_SLI;
				end else if (btnL == 1) begin
					next_state = S3_BOX;
				end else if (btnU == 1) begin
					next_state = S4_SPL;
				end */else begin
					next_state = S0_RESET;
				end
			end
			S1_MAP01: begin
				next_state = S1_MAP01;
			end
		endcase
	end
	
endmodule