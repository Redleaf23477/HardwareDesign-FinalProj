
/////////////////////////////////////////////////////////////////
// Constants Define
/////////////////////////////////////////////////////////////////

// player moving state

`define MOVE_STOP  3'd0
`define MOVE_DOWN  3'd1
`define MOVE_UP    3'd2
`define MOVE_LEFT  3'd3
`define MOVE_RIGHT 3'd4

// map size

`define MAP_ROW    10
`define MAP_COL    20

// map state

`define MAP_MAP0   3'd0
`define MAP_MAP1   3'd1

// shortest path state

`define STAT_STABLE 3'd0
`define STAT_INIT   3'd1
`define STAT_RELAX  3'd2


module bellman_ford_shortest_path(
	input clk,                         // faster clock
	input rst,
	input [9:0] player_r,
	input [9:0] player_c,
	
	input [2:0] map_stat,              // current map
	
	input [9:0] query_r0,
	input [9:0] query_c0,
	output [2:0] sp_dir0,               // shortest path backtrack on (query_r0, query_c0)
	output [9:0] sp_dist0,              // shortest path distance on (query_r0, query_c0)
	
	input [9:0] query_r1,
	input [9:0] query_c1,
	output [2:0] sp_dir1,
	output [9:0] sp_dist1,
	
	input [9:0] query_r2,
	input [9:0] query_c2,
	output [2:0] sp_dir2,
	output [9:0] sp_dist2,
	
	input [9:0] query_r3,
	input [9:0] query_c3,
	output [2:0] sp_dir3,
	output [9:0] sp_dist3,
	
	input [9:0] query_r4,
	input [9:0] query_c4,
	output [2:0] sp_dir4,
	output [9:0] sp_dist4
);

	reg [2:0] backtrack [0:9][0:19], nxt_backtrack[0:9][0:19];           // shortest path backtrack
	reg [9:0] shortest_dist [0:9][0:19], nxt_shortest_dist[0:9][0:19];   // shortest path distance

	// 0th query
	assign sp_dir0 = backtrack[query_r0][query_c0];
	assign sp_dist0 = shortest_dist[query_r0][query_c0];
	
	// 1st query
	assign sp_dir1 = backtrack[query_r1][query_c1];
	assign sp_dist1 = shortest_dist[query_r1][query_c1];
	
	// 2st query
	assign sp_dir2 = backtrack[query_r2][query_c2];
	assign sp_dist2 = shortest_dist[query_r2][query_c2];
	
	// 3st query
	assign sp_dir3 = backtrack[query_r3][query_c3];
	assign sp_dist3 = shortest_dist[query_r3][query_c3];
	
	// 4st query
	assign sp_dir4 = backtrack[query_r4][query_c4];
	assign sp_dist4 = shortest_dist[query_r4][query_c4];
	
	reg [9:0] prv_player_r, prv_player_c;
	reg [2:0] prv_map;
	reg [2:0] stat, nxt_stat;
	reg [9:0] loop_cnt, nxt_loop_cnt;

	// fsm with state
	always@(posedge clk, posedge rst) begin
		if(rst == 1'b1) begin
			stat <= `STAT_INIT;
			prv_player_r <= player_r;
			prv_player_c <= player_c;
			prv_map <= map_stat;
			loop_cnt <= 0;
		end else begin
			stat <= nxt_stat;
			prv_player_r <= player_r;
			prv_player_c <= player_c;
			prv_map <= map_stat;
			loop_cnt <= nxt_loop_cnt;
		end
	end
	always@(*) begin
		nxt_stat = stat;
		nxt_loop_cnt = loop_cnt;
		case(stat)
			`STAT_STABLE: begin
				if(map_stat == `MAP_MAP0 && (prv_player_r != player_r || prv_player_c != player_c )) begin
					nxt_stat = `STAT_INIT;
				end
			end
			`STAT_INIT: begin
				nxt_stat = `STAT_RELAX;
				nxt_loop_cnt = `MAP_ROW * `MAP_COL;
			end
			`STAT_RELAX: begin
				if(loop_cnt == 0) begin
					nxt_stat = `STAT_STABLE;
				end else begin
					nxt_loop_cnt = loop_cnt-1;
				end
			end
			default: begin
				nxt_stat = `STAT_STABLE;
				nxt_loop_cnt = 0;
			end
		endcase
	end
	
	// bellman ford relax
	always@(posedge clk) begin
		shift_backtrack;               // task
		shift_shortest_dist;           // task
	end
	always@(*) begin
		case(stat)
		`STAT_INIT: begin
			init_backtrack_map0;
			bf_init_shortest_path;
		end
		`STAT_RELAX: begin
			relax_backtrack_map0;
			relax_shortest_dist_map0;
		end
		default: begin
			shift_nxt_backtrack;           // task
			shift_nxt_shortest_dist;       // task
		end
		endcase
	end
	
	
	// tasks
task init_backtrack_map0;
begin
nxt_backtrack[0][0] <= `MOVE_STOP;
nxt_backtrack[0][1] <= `MOVE_STOP;
nxt_backtrack[0][2] <= `MOVE_STOP;
nxt_backtrack[0][3] <= `MOVE_STOP;
nxt_backtrack[0][4] <= `MOVE_STOP;
nxt_backtrack[0][5] <= `MOVE_STOP;
nxt_backtrack[0][6] <= `MOVE_STOP;
nxt_backtrack[0][7] <= `MOVE_STOP;
nxt_backtrack[0][8] <= `MOVE_STOP;
nxt_backtrack[0][9] <= `MOVE_STOP;
nxt_backtrack[0][10] <= `MOVE_STOP;
nxt_backtrack[0][11] <= `MOVE_STOP;
nxt_backtrack[0][12] <= `MOVE_STOP;
nxt_backtrack[0][13] <= `MOVE_STOP;
nxt_backtrack[0][14] <= `MOVE_STOP;
nxt_backtrack[0][15] <= `MOVE_STOP;
nxt_backtrack[0][16] <= `MOVE_STOP;
nxt_backtrack[0][17] <= `MOVE_STOP;
nxt_backtrack[0][18] <= `MOVE_STOP;
nxt_backtrack[0][19] <= `MOVE_STOP;
nxt_backtrack[1][0] <= `MOVE_STOP;
nxt_backtrack[1][1] <= `MOVE_RIGHT;
nxt_backtrack[1][2] <= `MOVE_RIGHT;
nxt_backtrack[1][3] <= `MOVE_DOWN;
nxt_backtrack[1][4] <= `MOVE_STOP;
nxt_backtrack[1][5] <= `MOVE_STOP;
nxt_backtrack[1][6] <= `MOVE_STOP;
nxt_backtrack[1][7] <= `MOVE_DOWN;
nxt_backtrack[1][8] <= `MOVE_STOP;
nxt_backtrack[1][9] <= `MOVE_STOP;
nxt_backtrack[1][10] <= `MOVE_DOWN;
nxt_backtrack[1][11] <= `MOVE_LEFT;
nxt_backtrack[1][12] <= `MOVE_LEFT;
nxt_backtrack[1][13] <= `MOVE_LEFT;
nxt_backtrack[1][14] <= `MOVE_LEFT;
nxt_backtrack[1][15] <= `MOVE_LEFT;
nxt_backtrack[1][16] <= `MOVE_LEFT;
nxt_backtrack[1][17] <= `MOVE_LEFT;
nxt_backtrack[1][18] <= `MOVE_DOWN;
nxt_backtrack[1][19] <= `MOVE_STOP;
nxt_backtrack[2][0] <= `MOVE_STOP;
nxt_backtrack[2][1] <= `MOVE_UP;
nxt_backtrack[2][2] <= `MOVE_STOP;
nxt_backtrack[2][3] <= `MOVE_DOWN;
nxt_backtrack[2][4] <= `MOVE_STOP;
nxt_backtrack[2][5] <= `MOVE_STOP;
nxt_backtrack[2][6] <= `MOVE_STOP;
nxt_backtrack[2][7] <= `MOVE_RIGHT;
nxt_backtrack[2][8] <= `MOVE_DOWN;
nxt_backtrack[2][9] <= `MOVE_LEFT;
nxt_backtrack[2][10] <= `MOVE_LEFT;
nxt_backtrack[2][11] <= `MOVE_STOP;
nxt_backtrack[2][12] <= `MOVE_STOP;
nxt_backtrack[2][13] <= `MOVE_STOP;
nxt_backtrack[2][14] <= `MOVE_UP;
nxt_backtrack[2][15] <= `MOVE_STOP;
nxt_backtrack[2][16] <= `MOVE_STOP;
nxt_backtrack[2][17] <= `MOVE_STOP;
nxt_backtrack[2][18] <= `MOVE_DOWN;
nxt_backtrack[2][19] <= `MOVE_STOP;
nxt_backtrack[3][0] <= `MOVE_STOP;
nxt_backtrack[3][1] <= `MOVE_UP;
nxt_backtrack[3][2] <= `MOVE_STOP;
nxt_backtrack[3][3] <= `MOVE_RIGHT;
nxt_backtrack[3][4] <= `MOVE_LEFT;
nxt_backtrack[3][5] <= `MOVE_LEFT;
nxt_backtrack[3][6] <= `MOVE_LEFT;
nxt_backtrack[3][7] <= `MOVE_STOP;
nxt_backtrack[3][8] <= `MOVE_DOWN;
nxt_backtrack[3][9] <= `MOVE_STOP;
nxt_backtrack[3][10] <= `MOVE_STOP;
nxt_backtrack[3][11] <= `MOVE_STOP;
nxt_backtrack[3][12] <= `MOVE_STOP;
nxt_backtrack[3][13] <= `MOVE_STOP;
nxt_backtrack[3][14] <= `MOVE_STOP;
nxt_backtrack[3][15] <= `MOVE_STOP;
nxt_backtrack[3][16] <= `MOVE_DOWN;
nxt_backtrack[3][17] <= `MOVE_LEFT;
nxt_backtrack[3][18] <= `MOVE_LEFT;
nxt_backtrack[3][19] <= `MOVE_STOP;
nxt_backtrack[4][0] <= `MOVE_STOP;
nxt_backtrack[4][1] <= `MOVE_UP;
nxt_backtrack[4][2] <= `MOVE_STOP;
nxt_backtrack[4][3] <= `MOVE_UP;
nxt_backtrack[4][4] <= `MOVE_STOP;
nxt_backtrack[4][5] <= `MOVE_UP;
nxt_backtrack[4][6] <= `MOVE_STOP;
nxt_backtrack[4][7] <= `MOVE_STOP;
nxt_backtrack[4][8] <= `MOVE_DOWN;
nxt_backtrack[4][9] <= `MOVE_STOP;
nxt_backtrack[4][10] <= `MOVE_STOP;
nxt_backtrack[4][11] <= `MOVE_STOP;
nxt_backtrack[4][12] <= `MOVE_STOP;
nxt_backtrack[4][13] <= `MOVE_DOWN;
nxt_backtrack[4][14] <= `MOVE_LEFT;
nxt_backtrack[4][15] <= `MOVE_LEFT;
nxt_backtrack[4][16] <= `MOVE_LEFT;
nxt_backtrack[4][17] <= `MOVE_STOP;
nxt_backtrack[4][18] <= `MOVE_STOP;
nxt_backtrack[4][19] <= `MOVE_STOP;
nxt_backtrack[5][0] <= `MOVE_STOP;
nxt_backtrack[5][1] <= `MOVE_STOP;
nxt_backtrack[5][2] <= `MOVE_STOP;
nxt_backtrack[5][3] <= `MOVE_STOP;
nxt_backtrack[5][4] <= `MOVE_STOP;
nxt_backtrack[5][5] <= `MOVE_UP;
nxt_backtrack[5][6] <= `MOVE_LEFT;
nxt_backtrack[5][7] <= `MOVE_LEFT;
nxt_backtrack[5][8] <= `MOVE_LEFT;
nxt_backtrack[5][9] <= `MOVE_LEFT;
nxt_backtrack[5][10] <= `MOVE_LEFT;
nxt_backtrack[5][11] <= `MOVE_LEFT;
nxt_backtrack[5][12] <= `MOVE_LEFT;
nxt_backtrack[5][13] <= `MOVE_LEFT;
nxt_backtrack[5][14] <= `MOVE_STOP;
nxt_backtrack[5][15] <= `MOVE_STOP;
nxt_backtrack[5][16] <= `MOVE_UP;
nxt_backtrack[5][17] <= `MOVE_LEFT;
nxt_backtrack[5][18] <= `MOVE_LEFT;
nxt_backtrack[5][19] <= `MOVE_STOP;
nxt_backtrack[6][0] <= `MOVE_STOP;
nxt_backtrack[6][1] <= `MOVE_DOWN;
nxt_backtrack[6][2] <= `MOVE_STOP;
nxt_backtrack[6][3] <= `MOVE_RIGHT;
nxt_backtrack[6][4] <= `MOVE_RIGHT;
nxt_backtrack[6][5] <= `MOVE_UP;
nxt_backtrack[6][6] <= `MOVE_UP;
nxt_backtrack[6][7] <= `MOVE_STOP;
nxt_backtrack[6][8] <= `MOVE_UP;
nxt_backtrack[6][9] <= `MOVE_STOP;
nxt_backtrack[6][10] <= `MOVE_STOP;
nxt_backtrack[6][11] <= `MOVE_STOP;
nxt_backtrack[6][12] <= `MOVE_STOP;
nxt_backtrack[6][13] <= `MOVE_UP;
nxt_backtrack[6][14] <= `MOVE_STOP;
nxt_backtrack[6][15] <= `MOVE_STOP;
nxt_backtrack[6][16] <= `MOVE_STOP;
nxt_backtrack[6][17] <= `MOVE_STOP;
nxt_backtrack[6][18] <= `MOVE_UP;
nxt_backtrack[6][19] <= `MOVE_STOP;
nxt_backtrack[7][0] <= `MOVE_STOP;
nxt_backtrack[7][1] <= `MOVE_DOWN;
nxt_backtrack[7][2] <= `MOVE_STOP;
nxt_backtrack[7][3] <= `MOVE_UP;
nxt_backtrack[7][4] <= `MOVE_STOP;
nxt_backtrack[7][5] <= `MOVE_STOP;
nxt_backtrack[7][6] <= `MOVE_UP;
nxt_backtrack[7][7] <= `MOVE_STOP;
nxt_backtrack[7][8] <= `MOVE_UP;
nxt_backtrack[7][9] <= `MOVE_LEFT;
nxt_backtrack[7][10] <= `MOVE_STOP;
nxt_backtrack[7][11] <= `MOVE_STOP;
nxt_backtrack[7][12] <= `MOVE_DOWN;
nxt_backtrack[7][13] <= `MOVE_UP;
nxt_backtrack[7][14] <= `MOVE_LEFT;
nxt_backtrack[7][15] <= `MOVE_LEFT;
nxt_backtrack[7][16] <= `MOVE_LEFT;
nxt_backtrack[7][17] <= `MOVE_STOP;
nxt_backtrack[7][18] <= `MOVE_DOWN;
nxt_backtrack[7][19] <= `MOVE_STOP;
nxt_backtrack[8][0] <= `MOVE_STOP;
nxt_backtrack[8][1] <= `MOVE_RIGHT;
nxt_backtrack[8][2] <= `MOVE_RIGHT;
nxt_backtrack[8][3] <= `MOVE_UP;
nxt_backtrack[8][4] <= `MOVE_STOP;
nxt_backtrack[8][5] <= `MOVE_STOP;
nxt_backtrack[8][6] <= `MOVE_UP;
nxt_backtrack[8][7] <= `MOVE_STOP;
nxt_backtrack[8][8] <= `MOVE_STOP;
nxt_backtrack[8][9] <= `MOVE_UP;
nxt_backtrack[8][10] <= `MOVE_LEFT;
nxt_backtrack[8][11] <= `MOVE_LEFT;
nxt_backtrack[8][12] <= `MOVE_LEFT;
nxt_backtrack[8][13] <= `MOVE_STOP;
nxt_backtrack[8][14] <= `MOVE_STOP;
nxt_backtrack[8][15] <= `MOVE_STOP;
nxt_backtrack[8][16] <= `MOVE_UP;
nxt_backtrack[8][17] <= `MOVE_LEFT;
nxt_backtrack[8][18] <= `MOVE_LEFT;
nxt_backtrack[8][19] <= `MOVE_STOP;
nxt_backtrack[9][0] <= `MOVE_STOP;
nxt_backtrack[9][1] <= `MOVE_STOP;
nxt_backtrack[9][2] <= `MOVE_STOP;
nxt_backtrack[9][3] <= `MOVE_STOP;
nxt_backtrack[9][4] <= `MOVE_STOP;
nxt_backtrack[9][5] <= `MOVE_STOP;
nxt_backtrack[9][6] <= `MOVE_STOP;
nxt_backtrack[9][7] <= `MOVE_STOP;
nxt_backtrack[9][8] <= `MOVE_STOP;
nxt_backtrack[9][9] <= `MOVE_STOP;
nxt_backtrack[9][10] <= `MOVE_STOP;
nxt_backtrack[9][11] <= `MOVE_STOP;
nxt_backtrack[9][12] <= `MOVE_STOP;
nxt_backtrack[9][13] <= `MOVE_STOP;
nxt_backtrack[9][14] <= `MOVE_STOP;
nxt_backtrack[9][15] <= `MOVE_STOP;
nxt_backtrack[9][16] <= `MOVE_STOP;
nxt_backtrack[9][17] <= `MOVE_STOP;
nxt_backtrack[9][18] <= `MOVE_STOP;
nxt_backtrack[9][19] <= `MOVE_STOP;
end
endtask
task relax_backtrack_map0;
begin
nxt_backtrack[0][0] <= backtrack[0][0];
nxt_backtrack[0][1] <= backtrack[0][1];
nxt_backtrack[0][2] <= backtrack[0][2];
nxt_backtrack[0][3] <= backtrack[0][3];
nxt_backtrack[0][4] <= backtrack[0][4];
nxt_backtrack[0][5] <= backtrack[0][5];
nxt_backtrack[0][6] <= backtrack[0][6];
nxt_backtrack[0][7] <= backtrack[0][7];
nxt_backtrack[0][8] <= backtrack[0][8];
nxt_backtrack[0][9] <= backtrack[0][9];
nxt_backtrack[0][10] <= backtrack[0][10];
nxt_backtrack[0][11] <= backtrack[0][11];
nxt_backtrack[0][12] <= backtrack[0][12];
nxt_backtrack[0][13] <= backtrack[0][13];
nxt_backtrack[0][14] <= backtrack[0][14];
nxt_backtrack[0][15] <= backtrack[0][15];
nxt_backtrack[0][16] <= backtrack[0][16];
nxt_backtrack[0][17] <= backtrack[0][17];
nxt_backtrack[0][18] <= backtrack[0][18];
nxt_backtrack[0][19] <= backtrack[0][19];
nxt_backtrack[1][0] <= backtrack[1][0];
nxt_backtrack[1][1] <= relax_dir(0,1,2,1,1,0,1,2,shortest_dist[1][1],backtrack[1][1]);
nxt_backtrack[1][2] <= relax_dir(0,2,2,2,1,1,1,3,shortest_dist[1][2],backtrack[1][2]);
nxt_backtrack[1][3] <= relax_dir(0,3,2,3,1,2,1,4,shortest_dist[1][3],backtrack[1][3]);
nxt_backtrack[1][4] <= backtrack[1][4];
nxt_backtrack[1][5] <= backtrack[1][5];
nxt_backtrack[1][6] <= backtrack[1][6];
nxt_backtrack[1][7] <= relax_dir(0,7,2,7,1,6,1,8,shortest_dist[1][7],backtrack[1][7]);
nxt_backtrack[1][8] <= backtrack[1][8];
nxt_backtrack[1][9] <= backtrack[1][9];
nxt_backtrack[1][10] <= relax_dir(0,10,2,10,1,9,1,11,shortest_dist[1][10],backtrack[1][10]);
nxt_backtrack[1][11] <= relax_dir(0,11,2,11,1,10,1,12,shortest_dist[1][11],backtrack[1][11]);
nxt_backtrack[1][12] <= relax_dir(0,12,2,12,1,11,1,13,shortest_dist[1][12],backtrack[1][12]);
nxt_backtrack[1][13] <= relax_dir(0,13,2,13,1,12,1,14,shortest_dist[1][13],backtrack[1][13]);
nxt_backtrack[1][14] <= relax_dir(0,14,2,14,1,13,1,15,shortest_dist[1][14],backtrack[1][14]);
nxt_backtrack[1][15] <= relax_dir(0,15,2,15,1,14,1,16,shortest_dist[1][15],backtrack[1][15]);
nxt_backtrack[1][16] <= relax_dir(0,16,2,16,1,15,1,17,shortest_dist[1][16],backtrack[1][16]);
nxt_backtrack[1][17] <= relax_dir(0,17,2,17,1,16,1,18,shortest_dist[1][17],backtrack[1][17]);
nxt_backtrack[1][18] <= relax_dir(0,18,2,18,1,17,1,19,shortest_dist[1][18],backtrack[1][18]);
nxt_backtrack[1][19] <= backtrack[1][19];
nxt_backtrack[2][0] <= backtrack[2][0];
nxt_backtrack[2][1] <= relax_dir(1,1,3,1,2,0,2,2,shortest_dist[2][1],backtrack[2][1]);
nxt_backtrack[2][2] <= backtrack[2][2];
nxt_backtrack[2][3] <= relax_dir(1,3,3,3,2,2,2,4,shortest_dist[2][3],backtrack[2][3]);
nxt_backtrack[2][4] <= backtrack[2][4];
nxt_backtrack[2][5] <= backtrack[2][5];
nxt_backtrack[2][6] <= backtrack[2][6];
nxt_backtrack[2][7] <= relax_dir(1,7,3,7,2,6,2,8,shortest_dist[2][7],backtrack[2][7]);
nxt_backtrack[2][8] <= relax_dir(1,8,3,8,2,7,2,9,shortest_dist[2][8],backtrack[2][8]);
nxt_backtrack[2][9] <= relax_dir(1,9,3,9,2,8,2,10,shortest_dist[2][9],backtrack[2][9]);
nxt_backtrack[2][10] <= relax_dir(1,10,3,10,2,9,2,11,shortest_dist[2][10],backtrack[2][10]);
nxt_backtrack[2][11] <= backtrack[2][11];
nxt_backtrack[2][12] <= backtrack[2][12];
nxt_backtrack[2][13] <= backtrack[2][13];
nxt_backtrack[2][14] <= relax_dir(1,14,3,14,2,13,2,15,shortest_dist[2][14],backtrack[2][14]);
nxt_backtrack[2][15] <= backtrack[2][15];
nxt_backtrack[2][16] <= backtrack[2][16];
nxt_backtrack[2][17] <= backtrack[2][17];
nxt_backtrack[2][18] <= relax_dir(1,18,3,18,2,17,2,19,shortest_dist[2][18],backtrack[2][18]);
nxt_backtrack[2][19] <= backtrack[2][19];
nxt_backtrack[3][0] <= backtrack[3][0];
nxt_backtrack[3][1] <= relax_dir(2,1,4,1,3,0,3,2,shortest_dist[3][1],backtrack[3][1]);
nxt_backtrack[3][2] <= backtrack[3][2];
nxt_backtrack[3][3] <= relax_dir(2,3,4,3,3,2,3,4,shortest_dist[3][3],backtrack[3][3]);
nxt_backtrack[3][4] <= relax_dir(2,4,4,4,3,3,3,5,shortest_dist[3][4],backtrack[3][4]);
nxt_backtrack[3][5] <= relax_dir(2,5,4,5,3,4,3,6,shortest_dist[3][5],backtrack[3][5]);
nxt_backtrack[3][6] <= relax_dir(2,6,4,6,3,5,3,7,shortest_dist[3][6],backtrack[3][6]);
nxt_backtrack[3][7] <= backtrack[3][7];
nxt_backtrack[3][8] <= relax_dir(2,8,4,8,3,7,3,9,shortest_dist[3][8],backtrack[3][8]);
nxt_backtrack[3][9] <= backtrack[3][9];
nxt_backtrack[3][10] <= backtrack[3][10];
nxt_backtrack[3][11] <= backtrack[3][11];
nxt_backtrack[3][12] <= backtrack[3][12];
nxt_backtrack[3][13] <= backtrack[3][13];
nxt_backtrack[3][14] <= backtrack[3][14];
nxt_backtrack[3][15] <= backtrack[3][15];
nxt_backtrack[3][16] <= relax_dir(2,16,4,16,3,15,3,17,shortest_dist[3][16],backtrack[3][16]);
nxt_backtrack[3][17] <= relax_dir(2,17,4,17,3,16,3,18,shortest_dist[3][17],backtrack[3][17]);
nxt_backtrack[3][18] <= relax_dir(2,18,4,18,3,17,3,19,shortest_dist[3][18],backtrack[3][18]);
nxt_backtrack[3][19] <= backtrack[3][19];
nxt_backtrack[4][0] <= backtrack[4][0];
nxt_backtrack[4][1] <= relax_dir(3,1,5,1,4,0,4,2,shortest_dist[4][1],backtrack[4][1]);
nxt_backtrack[4][2] <= backtrack[4][2];
nxt_backtrack[4][3] <= relax_dir(3,3,5,3,4,2,4,4,shortest_dist[4][3],backtrack[4][3]);
nxt_backtrack[4][4] <= backtrack[4][4];
nxt_backtrack[4][5] <= relax_dir(3,5,5,5,4,4,4,6,shortest_dist[4][5],backtrack[4][5]);
nxt_backtrack[4][6] <= backtrack[4][6];
nxt_backtrack[4][7] <= backtrack[4][7];
nxt_backtrack[4][8] <= relax_dir(3,8,5,8,4,7,4,9,shortest_dist[4][8],backtrack[4][8]);
nxt_backtrack[4][9] <= backtrack[4][9];
nxt_backtrack[4][10] <= backtrack[4][10];
nxt_backtrack[4][11] <= backtrack[4][11];
nxt_backtrack[4][12] <= backtrack[4][12];
nxt_backtrack[4][13] <= relax_dir(3,13,5,13,4,12,4,14,shortest_dist[4][13],backtrack[4][13]);
nxt_backtrack[4][14] <= relax_dir(3,14,5,14,4,13,4,15,shortest_dist[4][14],backtrack[4][14]);
nxt_backtrack[4][15] <= relax_dir(3,15,5,15,4,14,4,16,shortest_dist[4][15],backtrack[4][15]);
nxt_backtrack[4][16] <= relax_dir(3,16,5,16,4,15,4,17,shortest_dist[4][16],backtrack[4][16]);
nxt_backtrack[4][17] <= backtrack[4][17];
nxt_backtrack[4][18] <= backtrack[4][18];
nxt_backtrack[4][19] <= backtrack[4][19];
nxt_backtrack[5][0] <= backtrack[5][0];
nxt_backtrack[5][1] <= backtrack[5][1];
nxt_backtrack[5][2] <= backtrack[5][2];
nxt_backtrack[5][3] <= backtrack[5][3];
nxt_backtrack[5][4] <= backtrack[5][4];
nxt_backtrack[5][5] <= relax_dir(4,5,6,5,5,4,5,6,shortest_dist[5][5],backtrack[5][5]);
nxt_backtrack[5][6] <= relax_dir(4,6,6,6,5,5,5,7,shortest_dist[5][6],backtrack[5][6]);
nxt_backtrack[5][7] <= relax_dir(4,7,6,7,5,6,5,8,shortest_dist[5][7],backtrack[5][7]);
nxt_backtrack[5][8] <= relax_dir(4,8,6,8,5,7,5,9,shortest_dist[5][8],backtrack[5][8]);
nxt_backtrack[5][9] <= relax_dir(4,9,6,9,5,8,5,10,shortest_dist[5][9],backtrack[5][9]);
nxt_backtrack[5][10] <= relax_dir(4,10,6,10,5,9,5,11,shortest_dist[5][10],backtrack[5][10]);
nxt_backtrack[5][11] <= relax_dir(4,11,6,11,5,10,5,12,shortest_dist[5][11],backtrack[5][11]);
nxt_backtrack[5][12] <= relax_dir(4,12,6,12,5,11,5,13,shortest_dist[5][12],backtrack[5][12]);
nxt_backtrack[5][13] <= relax_dir(4,13,6,13,5,12,5,14,shortest_dist[5][13],backtrack[5][13]);
nxt_backtrack[5][14] <= backtrack[5][14];
nxt_backtrack[5][15] <= backtrack[5][15];
nxt_backtrack[5][16] <= relax_dir(4,16,6,16,5,15,5,17,shortest_dist[5][16],backtrack[5][16]);
nxt_backtrack[5][17] <= relax_dir(4,17,6,17,5,16,5,18,shortest_dist[5][17],backtrack[5][17]);
nxt_backtrack[5][18] <= relax_dir(4,18,6,18,5,17,5,19,shortest_dist[5][18],backtrack[5][18]);
nxt_backtrack[5][19] <= backtrack[5][19];
nxt_backtrack[6][0] <= backtrack[6][0];
nxt_backtrack[6][1] <= relax_dir(5,1,7,1,6,0,6,2,shortest_dist[6][1],backtrack[6][1]);
nxt_backtrack[6][2] <= backtrack[6][2];
nxt_backtrack[6][3] <= relax_dir(5,3,7,3,6,2,6,4,shortest_dist[6][3],backtrack[6][3]);
nxt_backtrack[6][4] <= relax_dir(5,4,7,4,6,3,6,5,shortest_dist[6][4],backtrack[6][4]);
nxt_backtrack[6][5] <= relax_dir(5,5,7,5,6,4,6,6,shortest_dist[6][5],backtrack[6][5]);
nxt_backtrack[6][6] <= relax_dir(5,6,7,6,6,5,6,7,shortest_dist[6][6],backtrack[6][6]);
nxt_backtrack[6][7] <= backtrack[6][7];
nxt_backtrack[6][8] <= relax_dir(5,8,7,8,6,7,6,9,shortest_dist[6][8],backtrack[6][8]);
nxt_backtrack[6][9] <= backtrack[6][9];
nxt_backtrack[6][10] <= backtrack[6][10];
nxt_backtrack[6][11] <= backtrack[6][11];
nxt_backtrack[6][12] <= backtrack[6][12];
nxt_backtrack[6][13] <= relax_dir(5,13,7,13,6,12,6,14,shortest_dist[6][13],backtrack[6][13]);
nxt_backtrack[6][14] <= backtrack[6][14];
nxt_backtrack[6][15] <= backtrack[6][15];
nxt_backtrack[6][16] <= backtrack[6][16];
nxt_backtrack[6][17] <= backtrack[6][17];
nxt_backtrack[6][18] <= relax_dir(5,18,7,18,6,17,6,19,shortest_dist[6][18],backtrack[6][18]);
nxt_backtrack[6][19] <= backtrack[6][19];
nxt_backtrack[7][0] <= backtrack[7][0];
nxt_backtrack[7][1] <= relax_dir(6,1,8,1,7,0,7,2,shortest_dist[7][1],backtrack[7][1]);
nxt_backtrack[7][2] <= backtrack[7][2];
nxt_backtrack[7][3] <= relax_dir(6,3,8,3,7,2,7,4,shortest_dist[7][3],backtrack[7][3]);
nxt_backtrack[7][4] <= backtrack[7][4];
nxt_backtrack[7][5] <= backtrack[7][5];
nxt_backtrack[7][6] <= relax_dir(6,6,8,6,7,5,7,7,shortest_dist[7][6],backtrack[7][6]);
nxt_backtrack[7][7] <= backtrack[7][7];
nxt_backtrack[7][8] <= relax_dir(6,8,8,8,7,7,7,9,shortest_dist[7][8],backtrack[7][8]);
nxt_backtrack[7][9] <= relax_dir(6,9,8,9,7,8,7,10,shortest_dist[7][9],backtrack[7][9]);
nxt_backtrack[7][10] <= backtrack[7][10];
nxt_backtrack[7][11] <= backtrack[7][11];
nxt_backtrack[7][12] <= relax_dir(6,12,8,12,7,11,7,13,shortest_dist[7][12],backtrack[7][12]);
nxt_backtrack[7][13] <= relax_dir(6,13,8,13,7,12,7,14,shortest_dist[7][13],backtrack[7][13]);
nxt_backtrack[7][14] <= relax_dir(6,14,8,14,7,13,7,15,shortest_dist[7][14],backtrack[7][14]);
nxt_backtrack[7][15] <= relax_dir(6,15,8,15,7,14,7,16,shortest_dist[7][15],backtrack[7][15]);
nxt_backtrack[7][16] <= relax_dir(6,16,8,16,7,15,7,17,shortest_dist[7][16],backtrack[7][16]);
nxt_backtrack[7][17] <= backtrack[7][17];
nxt_backtrack[7][18] <= relax_dir(6,18,8,18,7,17,7,19,shortest_dist[7][18],backtrack[7][18]);
nxt_backtrack[7][19] <= backtrack[7][19];
nxt_backtrack[8][0] <= backtrack[8][0];
nxt_backtrack[8][1] <= relax_dir(7,1,9,1,8,0,8,2,shortest_dist[8][1],backtrack[8][1]);
nxt_backtrack[8][2] <= relax_dir(7,2,9,2,8,1,8,3,shortest_dist[8][2],backtrack[8][2]);
nxt_backtrack[8][3] <= relax_dir(7,3,9,3,8,2,8,4,shortest_dist[8][3],backtrack[8][3]);
nxt_backtrack[8][4] <= backtrack[8][4];
nxt_backtrack[8][5] <= backtrack[8][5];
nxt_backtrack[8][6] <= relax_dir(7,6,9,6,8,5,8,7,shortest_dist[8][6],backtrack[8][6]);
nxt_backtrack[8][7] <= backtrack[8][7];
nxt_backtrack[8][8] <= backtrack[8][8];
nxt_backtrack[8][9] <= relax_dir(7,9,9,9,8,8,8,10,shortest_dist[8][9],backtrack[8][9]);
nxt_backtrack[8][10] <= relax_dir(7,10,9,10,8,9,8,11,shortest_dist[8][10],backtrack[8][10]);
nxt_backtrack[8][11] <= relax_dir(7,11,9,11,8,10,8,12,shortest_dist[8][11],backtrack[8][11]);
nxt_backtrack[8][12] <= relax_dir(7,12,9,12,8,11,8,13,shortest_dist[8][12],backtrack[8][12]);
nxt_backtrack[8][13] <= backtrack[8][13];
nxt_backtrack[8][14] <= backtrack[8][14];
nxt_backtrack[8][15] <= backtrack[8][15];
nxt_backtrack[8][16] <= relax_dir(7,16,9,16,8,15,8,17,shortest_dist[8][16],backtrack[8][16]);
nxt_backtrack[8][17] <= relax_dir(7,17,9,17,8,16,8,18,shortest_dist[8][17],backtrack[8][17]);
nxt_backtrack[8][18] <= relax_dir(7,18,9,18,8,17,8,19,shortest_dist[8][18],backtrack[8][18]);
nxt_backtrack[8][19] <= backtrack[8][19];
nxt_backtrack[9][0] <= backtrack[9][0];
nxt_backtrack[9][1] <= backtrack[9][1];
nxt_backtrack[9][2] <= backtrack[9][2];
nxt_backtrack[9][3] <= backtrack[9][3];
nxt_backtrack[9][4] <= backtrack[9][4];
nxt_backtrack[9][5] <= backtrack[9][5];
nxt_backtrack[9][6] <= backtrack[9][6];
nxt_backtrack[9][7] <= backtrack[9][7];
nxt_backtrack[9][8] <= backtrack[9][8];
nxt_backtrack[9][9] <= backtrack[9][9];
nxt_backtrack[9][10] <= backtrack[9][10];
nxt_backtrack[9][11] <= backtrack[9][11];
nxt_backtrack[9][12] <= backtrack[9][12];
nxt_backtrack[9][13] <= backtrack[9][13];
nxt_backtrack[9][14] <= backtrack[9][14];
nxt_backtrack[9][15] <= backtrack[9][15];
nxt_backtrack[9][16] <= backtrack[9][16];
nxt_backtrack[9][17] <= backtrack[9][17];
nxt_backtrack[9][18] <= backtrack[9][18];
nxt_backtrack[9][19] <= backtrack[9][19];
end
endtask
task relax_shortest_dist_map0;
begin
nxt_shortest_dist[0][0] <= shortest_dist[0][0];
nxt_shortest_dist[0][1] <= shortest_dist[0][1];
nxt_shortest_dist[0][2] <= shortest_dist[0][2];
nxt_shortest_dist[0][3] <= shortest_dist[0][3];
nxt_shortest_dist[0][4] <= shortest_dist[0][4];
nxt_shortest_dist[0][5] <= shortest_dist[0][5];
nxt_shortest_dist[0][6] <= shortest_dist[0][6];
nxt_shortest_dist[0][7] <= shortest_dist[0][7];
nxt_shortest_dist[0][8] <= shortest_dist[0][8];
nxt_shortest_dist[0][9] <= shortest_dist[0][9];
nxt_shortest_dist[0][10] <= shortest_dist[0][10];
nxt_shortest_dist[0][11] <= shortest_dist[0][11];
nxt_shortest_dist[0][12] <= shortest_dist[0][12];
nxt_shortest_dist[0][13] <= shortest_dist[0][13];
nxt_shortest_dist[0][14] <= shortest_dist[0][14];
nxt_shortest_dist[0][15] <= shortest_dist[0][15];
nxt_shortest_dist[0][16] <= shortest_dist[0][16];
nxt_shortest_dist[0][17] <= shortest_dist[0][17];
nxt_shortest_dist[0][18] <= shortest_dist[0][18];
nxt_shortest_dist[0][19] <= shortest_dist[0][19];
nxt_shortest_dist[1][0] <= shortest_dist[1][0];
nxt_shortest_dist[1][1] <= relax_dist(0,1,2,1,1,0,1,2,shortest_dist[1][1]);
nxt_shortest_dist[1][2] <= relax_dist(0,2,2,2,1,1,1,3,shortest_dist[1][2]);
nxt_shortest_dist[1][3] <= relax_dist(0,3,2,3,1,2,1,4,shortest_dist[1][3]);
nxt_shortest_dist[1][4] <= shortest_dist[1][4];
nxt_shortest_dist[1][5] <= shortest_dist[1][5];
nxt_shortest_dist[1][6] <= shortest_dist[1][6];
nxt_shortest_dist[1][7] <= relax_dist(0,7,2,7,1,6,1,8,shortest_dist[1][7]);
nxt_shortest_dist[1][8] <= shortest_dist[1][8];
nxt_shortest_dist[1][9] <= shortest_dist[1][9];
nxt_shortest_dist[1][10] <= relax_dist(0,10,2,10,1,9,1,11,shortest_dist[1][10]);
nxt_shortest_dist[1][11] <= relax_dist(0,11,2,11,1,10,1,12,shortest_dist[1][11]);
nxt_shortest_dist[1][12] <= relax_dist(0,12,2,12,1,11,1,13,shortest_dist[1][12]);
nxt_shortest_dist[1][13] <= relax_dist(0,13,2,13,1,12,1,14,shortest_dist[1][13]);
nxt_shortest_dist[1][14] <= relax_dist(0,14,2,14,1,13,1,15,shortest_dist[1][14]);
nxt_shortest_dist[1][15] <= relax_dist(0,15,2,15,1,14,1,16,shortest_dist[1][15]);
nxt_shortest_dist[1][16] <= relax_dist(0,16,2,16,1,15,1,17,shortest_dist[1][16]);
nxt_shortest_dist[1][17] <= relax_dist(0,17,2,17,1,16,1,18,shortest_dist[1][17]);
nxt_shortest_dist[1][18] <= relax_dist(0,18,2,18,1,17,1,19,shortest_dist[1][18]);
nxt_shortest_dist[1][19] <= shortest_dist[1][19];
nxt_shortest_dist[2][0] <= shortest_dist[2][0];
nxt_shortest_dist[2][1] <= relax_dist(1,1,3,1,2,0,2,2,shortest_dist[2][1]);
nxt_shortest_dist[2][2] <= shortest_dist[2][2];
nxt_shortest_dist[2][3] <= relax_dist(1,3,3,3,2,2,2,4,shortest_dist[2][3]);
nxt_shortest_dist[2][4] <= shortest_dist[2][4];
nxt_shortest_dist[2][5] <= shortest_dist[2][5];
nxt_shortest_dist[2][6] <= shortest_dist[2][6];
nxt_shortest_dist[2][7] <= relax_dist(1,7,3,7,2,6,2,8,shortest_dist[2][7]);
nxt_shortest_dist[2][8] <= relax_dist(1,8,3,8,2,7,2,9,shortest_dist[2][8]);
nxt_shortest_dist[2][9] <= relax_dist(1,9,3,9,2,8,2,10,shortest_dist[2][9]);
nxt_shortest_dist[2][10] <= relax_dist(1,10,3,10,2,9,2,11,shortest_dist[2][10]);
nxt_shortest_dist[2][11] <= shortest_dist[2][11];
nxt_shortest_dist[2][12] <= shortest_dist[2][12];
nxt_shortest_dist[2][13] <= shortest_dist[2][13];
nxt_shortest_dist[2][14] <= relax_dist(1,14,3,14,2,13,2,15,shortest_dist[2][14]);
nxt_shortest_dist[2][15] <= shortest_dist[2][15];
nxt_shortest_dist[2][16] <= shortest_dist[2][16];
nxt_shortest_dist[2][17] <= shortest_dist[2][17];
nxt_shortest_dist[2][18] <= relax_dist(1,18,3,18,2,17,2,19,shortest_dist[2][18]);
nxt_shortest_dist[2][19] <= shortest_dist[2][19];
nxt_shortest_dist[3][0] <= shortest_dist[3][0];
nxt_shortest_dist[3][1] <= relax_dist(2,1,4,1,3,0,3,2,shortest_dist[3][1]);
nxt_shortest_dist[3][2] <= shortest_dist[3][2];
nxt_shortest_dist[3][3] <= relax_dist(2,3,4,3,3,2,3,4,shortest_dist[3][3]);
nxt_shortest_dist[3][4] <= relax_dist(2,4,4,4,3,3,3,5,shortest_dist[3][4]);
nxt_shortest_dist[3][5] <= relax_dist(2,5,4,5,3,4,3,6,shortest_dist[3][5]);
nxt_shortest_dist[3][6] <= relax_dist(2,6,4,6,3,5,3,7,shortest_dist[3][6]);
nxt_shortest_dist[3][7] <= shortest_dist[3][7];
nxt_shortest_dist[3][8] <= relax_dist(2,8,4,8,3,7,3,9,shortest_dist[3][8]);
nxt_shortest_dist[3][9] <= shortest_dist[3][9];
nxt_shortest_dist[3][10] <= shortest_dist[3][10];
nxt_shortest_dist[3][11] <= shortest_dist[3][11];
nxt_shortest_dist[3][12] <= shortest_dist[3][12];
nxt_shortest_dist[3][13] <= shortest_dist[3][13];
nxt_shortest_dist[3][14] <= shortest_dist[3][14];
nxt_shortest_dist[3][15] <= shortest_dist[3][15];
nxt_shortest_dist[3][16] <= relax_dist(2,16,4,16,3,15,3,17,shortest_dist[3][16]);
nxt_shortest_dist[3][17] <= relax_dist(2,17,4,17,3,16,3,18,shortest_dist[3][17]);
nxt_shortest_dist[3][18] <= relax_dist(2,18,4,18,3,17,3,19,shortest_dist[3][18]);
nxt_shortest_dist[3][19] <= shortest_dist[3][19];
nxt_shortest_dist[4][0] <= shortest_dist[4][0];
nxt_shortest_dist[4][1] <= relax_dist(3,1,5,1,4,0,4,2,shortest_dist[4][1]);
nxt_shortest_dist[4][2] <= shortest_dist[4][2];
nxt_shortest_dist[4][3] <= relax_dist(3,3,5,3,4,2,4,4,shortest_dist[4][3]);
nxt_shortest_dist[4][4] <= shortest_dist[4][4];
nxt_shortest_dist[4][5] <= relax_dist(3,5,5,5,4,4,4,6,shortest_dist[4][5]);
nxt_shortest_dist[4][6] <= shortest_dist[4][6];
nxt_shortest_dist[4][7] <= shortest_dist[4][7];
nxt_shortest_dist[4][8] <= relax_dist(3,8,5,8,4,7,4,9,shortest_dist[4][8]);
nxt_shortest_dist[4][9] <= shortest_dist[4][9];
nxt_shortest_dist[4][10] <= shortest_dist[4][10];
nxt_shortest_dist[4][11] <= shortest_dist[4][11];
nxt_shortest_dist[4][12] <= shortest_dist[4][12];
nxt_shortest_dist[4][13] <= relax_dist(3,13,5,13,4,12,4,14,shortest_dist[4][13]);
nxt_shortest_dist[4][14] <= relax_dist(3,14,5,14,4,13,4,15,shortest_dist[4][14]);
nxt_shortest_dist[4][15] <= relax_dist(3,15,5,15,4,14,4,16,shortest_dist[4][15]);
nxt_shortest_dist[4][16] <= relax_dist(3,16,5,16,4,15,4,17,shortest_dist[4][16]);
nxt_shortest_dist[4][17] <= shortest_dist[4][17];
nxt_shortest_dist[4][18] <= shortest_dist[4][18];
nxt_shortest_dist[4][19] <= shortest_dist[4][19];
nxt_shortest_dist[5][0] <= shortest_dist[5][0];
nxt_shortest_dist[5][1] <= shortest_dist[5][1];
nxt_shortest_dist[5][2] <= shortest_dist[5][2];
nxt_shortest_dist[5][3] <= shortest_dist[5][3];
nxt_shortest_dist[5][4] <= shortest_dist[5][4];
nxt_shortest_dist[5][5] <= relax_dist(4,5,6,5,5,4,5,6,shortest_dist[5][5]);
nxt_shortest_dist[5][6] <= relax_dist(4,6,6,6,5,5,5,7,shortest_dist[5][6]);
nxt_shortest_dist[5][7] <= relax_dist(4,7,6,7,5,6,5,8,shortest_dist[5][7]);
nxt_shortest_dist[5][8] <= relax_dist(4,8,6,8,5,7,5,9,shortest_dist[5][8]);
nxt_shortest_dist[5][9] <= relax_dist(4,9,6,9,5,8,5,10,shortest_dist[5][9]);
nxt_shortest_dist[5][10] <= relax_dist(4,10,6,10,5,9,5,11,shortest_dist[5][10]);
nxt_shortest_dist[5][11] <= relax_dist(4,11,6,11,5,10,5,12,shortest_dist[5][11]);
nxt_shortest_dist[5][12] <= relax_dist(4,12,6,12,5,11,5,13,shortest_dist[5][12]);
nxt_shortest_dist[5][13] <= relax_dist(4,13,6,13,5,12,5,14,shortest_dist[5][13]);
nxt_shortest_dist[5][14] <= shortest_dist[5][14];
nxt_shortest_dist[5][15] <= shortest_dist[5][15];
nxt_shortest_dist[5][16] <= relax_dist(4,16,6,16,5,15,5,17,shortest_dist[5][16]);
nxt_shortest_dist[5][17] <= relax_dist(4,17,6,17,5,16,5,18,shortest_dist[5][17]);
nxt_shortest_dist[5][18] <= relax_dist(4,18,6,18,5,17,5,19,shortest_dist[5][18]);
nxt_shortest_dist[5][19] <= shortest_dist[5][19];
nxt_shortest_dist[6][0] <= shortest_dist[6][0];
nxt_shortest_dist[6][1] <= relax_dist(5,1,7,1,6,0,6,2,shortest_dist[6][1]);
nxt_shortest_dist[6][2] <= shortest_dist[6][2];
nxt_shortest_dist[6][3] <= relax_dist(5,3,7,3,6,2,6,4,shortest_dist[6][3]);
nxt_shortest_dist[6][4] <= relax_dist(5,4,7,4,6,3,6,5,shortest_dist[6][4]);
nxt_shortest_dist[6][5] <= relax_dist(5,5,7,5,6,4,6,6,shortest_dist[6][5]);
nxt_shortest_dist[6][6] <= relax_dist(5,6,7,6,6,5,6,7,shortest_dist[6][6]);
nxt_shortest_dist[6][7] <= shortest_dist[6][7];
nxt_shortest_dist[6][8] <= relax_dist(5,8,7,8,6,7,6,9,shortest_dist[6][8]);
nxt_shortest_dist[6][9] <= shortest_dist[6][9];
nxt_shortest_dist[6][10] <= shortest_dist[6][10];
nxt_shortest_dist[6][11] <= shortest_dist[6][11];
nxt_shortest_dist[6][12] <= shortest_dist[6][12];
nxt_shortest_dist[6][13] <= relax_dist(5,13,7,13,6,12,6,14,shortest_dist[6][13]);
nxt_shortest_dist[6][14] <= shortest_dist[6][14];
nxt_shortest_dist[6][15] <= shortest_dist[6][15];
nxt_shortest_dist[6][16] <= shortest_dist[6][16];
nxt_shortest_dist[6][17] <= shortest_dist[6][17];
nxt_shortest_dist[6][18] <= relax_dist(5,18,7,18,6,17,6,19,shortest_dist[6][18]);
nxt_shortest_dist[6][19] <= shortest_dist[6][19];
nxt_shortest_dist[7][0] <= shortest_dist[7][0];
nxt_shortest_dist[7][1] <= relax_dist(6,1,8,1,7,0,7,2,shortest_dist[7][1]);
nxt_shortest_dist[7][2] <= shortest_dist[7][2];
nxt_shortest_dist[7][3] <= relax_dist(6,3,8,3,7,2,7,4,shortest_dist[7][3]);
nxt_shortest_dist[7][4] <= shortest_dist[7][4];
nxt_shortest_dist[7][5] <= shortest_dist[7][5];
nxt_shortest_dist[7][6] <= relax_dist(6,6,8,6,7,5,7,7,shortest_dist[7][6]);
nxt_shortest_dist[7][7] <= shortest_dist[7][7];
nxt_shortest_dist[7][8] <= relax_dist(6,8,8,8,7,7,7,9,shortest_dist[7][8]);
nxt_shortest_dist[7][9] <= relax_dist(6,9,8,9,7,8,7,10,shortest_dist[7][9]);
nxt_shortest_dist[7][10] <= shortest_dist[7][10];
nxt_shortest_dist[7][11] <= shortest_dist[7][11];
nxt_shortest_dist[7][12] <= relax_dist(6,12,8,12,7,11,7,13,shortest_dist[7][12]);
nxt_shortest_dist[7][13] <= relax_dist(6,13,8,13,7,12,7,14,shortest_dist[7][13]);
nxt_shortest_dist[7][14] <= relax_dist(6,14,8,14,7,13,7,15,shortest_dist[7][14]);
nxt_shortest_dist[7][15] <= relax_dist(6,15,8,15,7,14,7,16,shortest_dist[7][15]);
nxt_shortest_dist[7][16] <= relax_dist(6,16,8,16,7,15,7,17,shortest_dist[7][16]);
nxt_shortest_dist[7][17] <= shortest_dist[7][17];
nxt_shortest_dist[7][18] <= relax_dist(6,18,8,18,7,17,7,19,shortest_dist[7][18]);
nxt_shortest_dist[7][19] <= shortest_dist[7][19];
nxt_shortest_dist[8][0] <= shortest_dist[8][0];
nxt_shortest_dist[8][1] <= relax_dist(7,1,9,1,8,0,8,2,shortest_dist[8][1]);
nxt_shortest_dist[8][2] <= relax_dist(7,2,9,2,8,1,8,3,shortest_dist[8][2]);
nxt_shortest_dist[8][3] <= relax_dist(7,3,9,3,8,2,8,4,shortest_dist[8][3]);
nxt_shortest_dist[8][4] <= shortest_dist[8][4];
nxt_shortest_dist[8][5] <= shortest_dist[8][5];
nxt_shortest_dist[8][6] <= relax_dist(7,6,9,6,8,5,8,7,shortest_dist[8][6]);
nxt_shortest_dist[8][7] <= shortest_dist[8][7];
nxt_shortest_dist[8][8] <= shortest_dist[8][8];
nxt_shortest_dist[8][9] <= relax_dist(7,9,9,9,8,8,8,10,shortest_dist[8][9]);
nxt_shortest_dist[8][10] <= relax_dist(7,10,9,10,8,9,8,11,shortest_dist[8][10]);
nxt_shortest_dist[8][11] <= relax_dist(7,11,9,11,8,10,8,12,shortest_dist[8][11]);
nxt_shortest_dist[8][12] <= relax_dist(7,12,9,12,8,11,8,13,shortest_dist[8][12]);
nxt_shortest_dist[8][13] <= shortest_dist[8][13];
nxt_shortest_dist[8][14] <= shortest_dist[8][14];
nxt_shortest_dist[8][15] <= shortest_dist[8][15];
nxt_shortest_dist[8][16] <= relax_dist(7,16,9,16,8,15,8,17,shortest_dist[8][16]);
nxt_shortest_dist[8][17] <= relax_dist(7,17,9,17,8,16,8,18,shortest_dist[8][17]);
nxt_shortest_dist[8][18] <= relax_dist(7,18,9,18,8,17,8,19,shortest_dist[8][18]);
nxt_shortest_dist[8][19] <= shortest_dist[8][19];
nxt_shortest_dist[9][0] <= shortest_dist[9][0];
nxt_shortest_dist[9][1] <= shortest_dist[9][1];
nxt_shortest_dist[9][2] <= shortest_dist[9][2];
nxt_shortest_dist[9][3] <= shortest_dist[9][3];
nxt_shortest_dist[9][4] <= shortest_dist[9][4];
nxt_shortest_dist[9][5] <= shortest_dist[9][5];
nxt_shortest_dist[9][6] <= shortest_dist[9][6];
nxt_shortest_dist[9][7] <= shortest_dist[9][7];
nxt_shortest_dist[9][8] <= shortest_dist[9][8];
nxt_shortest_dist[9][9] <= shortest_dist[9][9];
nxt_shortest_dist[9][10] <= shortest_dist[9][10];
nxt_shortest_dist[9][11] <= shortest_dist[9][11];
nxt_shortest_dist[9][12] <= shortest_dist[9][12];
nxt_shortest_dist[9][13] <= shortest_dist[9][13];
nxt_shortest_dist[9][14] <= shortest_dist[9][14];
nxt_shortest_dist[9][15] <= shortest_dist[9][15];
nxt_shortest_dist[9][16] <= shortest_dist[9][16];
nxt_shortest_dist[9][17] <= shortest_dist[9][17];
nxt_shortest_dist[9][18] <= shortest_dist[9][18];
nxt_shortest_dist[9][19] <= shortest_dist[9][19];
end
endtask

task shift_backtrack;
begin
backtrack[0][0] <= nxt_backtrack[0][0];
backtrack[0][1] <= nxt_backtrack[0][1];
backtrack[0][2] <= nxt_backtrack[0][2];
backtrack[0][3] <= nxt_backtrack[0][3];
backtrack[0][4] <= nxt_backtrack[0][4];
backtrack[0][5] <= nxt_backtrack[0][5];
backtrack[0][6] <= nxt_backtrack[0][6];
backtrack[0][7] <= nxt_backtrack[0][7];
backtrack[0][8] <= nxt_backtrack[0][8];
backtrack[0][9] <= nxt_backtrack[0][9];
backtrack[0][10] <= nxt_backtrack[0][10];
backtrack[0][11] <= nxt_backtrack[0][11];
backtrack[0][12] <= nxt_backtrack[0][12];
backtrack[0][13] <= nxt_backtrack[0][13];
backtrack[0][14] <= nxt_backtrack[0][14];
backtrack[0][15] <= nxt_backtrack[0][15];
backtrack[0][16] <= nxt_backtrack[0][16];
backtrack[0][17] <= nxt_backtrack[0][17];
backtrack[0][18] <= nxt_backtrack[0][18];
backtrack[0][19] <= nxt_backtrack[0][19];
backtrack[1][0] <= nxt_backtrack[1][0];
backtrack[1][1] <= nxt_backtrack[1][1];
backtrack[1][2] <= nxt_backtrack[1][2];
backtrack[1][3] <= nxt_backtrack[1][3];
backtrack[1][4] <= nxt_backtrack[1][4];
backtrack[1][5] <= nxt_backtrack[1][5];
backtrack[1][6] <= nxt_backtrack[1][6];
backtrack[1][7] <= nxt_backtrack[1][7];
backtrack[1][8] <= nxt_backtrack[1][8];
backtrack[1][9] <= nxt_backtrack[1][9];
backtrack[1][10] <= nxt_backtrack[1][10];
backtrack[1][11] <= nxt_backtrack[1][11];
backtrack[1][12] <= nxt_backtrack[1][12];
backtrack[1][13] <= nxt_backtrack[1][13];
backtrack[1][14] <= nxt_backtrack[1][14];
backtrack[1][15] <= nxt_backtrack[1][15];
backtrack[1][16] <= nxt_backtrack[1][16];
backtrack[1][17] <= nxt_backtrack[1][17];
backtrack[1][18] <= nxt_backtrack[1][18];
backtrack[1][19] <= nxt_backtrack[1][19];
backtrack[2][0] <= nxt_backtrack[2][0];
backtrack[2][1] <= nxt_backtrack[2][1];
backtrack[2][2] <= nxt_backtrack[2][2];
backtrack[2][3] <= nxt_backtrack[2][3];
backtrack[2][4] <= nxt_backtrack[2][4];
backtrack[2][5] <= nxt_backtrack[2][5];
backtrack[2][6] <= nxt_backtrack[2][6];
backtrack[2][7] <= nxt_backtrack[2][7];
backtrack[2][8] <= nxt_backtrack[2][8];
backtrack[2][9] <= nxt_backtrack[2][9];
backtrack[2][10] <= nxt_backtrack[2][10];
backtrack[2][11] <= nxt_backtrack[2][11];
backtrack[2][12] <= nxt_backtrack[2][12];
backtrack[2][13] <= nxt_backtrack[2][13];
backtrack[2][14] <= nxt_backtrack[2][14];
backtrack[2][15] <= nxt_backtrack[2][15];
backtrack[2][16] <= nxt_backtrack[2][16];
backtrack[2][17] <= nxt_backtrack[2][17];
backtrack[2][18] <= nxt_backtrack[2][18];
backtrack[2][19] <= nxt_backtrack[2][19];
backtrack[3][0] <= nxt_backtrack[3][0];
backtrack[3][1] <= nxt_backtrack[3][1];
backtrack[3][2] <= nxt_backtrack[3][2];
backtrack[3][3] <= nxt_backtrack[3][3];
backtrack[3][4] <= nxt_backtrack[3][4];
backtrack[3][5] <= nxt_backtrack[3][5];
backtrack[3][6] <= nxt_backtrack[3][6];
backtrack[3][7] <= nxt_backtrack[3][7];
backtrack[3][8] <= nxt_backtrack[3][8];
backtrack[3][9] <= nxt_backtrack[3][9];
backtrack[3][10] <= nxt_backtrack[3][10];
backtrack[3][11] <= nxt_backtrack[3][11];
backtrack[3][12] <= nxt_backtrack[3][12];
backtrack[3][13] <= nxt_backtrack[3][13];
backtrack[3][14] <= nxt_backtrack[3][14];
backtrack[3][15] <= nxt_backtrack[3][15];
backtrack[3][16] <= nxt_backtrack[3][16];
backtrack[3][17] <= nxt_backtrack[3][17];
backtrack[3][18] <= nxt_backtrack[3][18];
backtrack[3][19] <= nxt_backtrack[3][19];
backtrack[4][0] <= nxt_backtrack[4][0];
backtrack[4][1] <= nxt_backtrack[4][1];
backtrack[4][2] <= nxt_backtrack[4][2];
backtrack[4][3] <= nxt_backtrack[4][3];
backtrack[4][4] <= nxt_backtrack[4][4];
backtrack[4][5] <= nxt_backtrack[4][5];
backtrack[4][6] <= nxt_backtrack[4][6];
backtrack[4][7] <= nxt_backtrack[4][7];
backtrack[4][8] <= nxt_backtrack[4][8];
backtrack[4][9] <= nxt_backtrack[4][9];
backtrack[4][10] <= nxt_backtrack[4][10];
backtrack[4][11] <= nxt_backtrack[4][11];
backtrack[4][12] <= nxt_backtrack[4][12];
backtrack[4][13] <= nxt_backtrack[4][13];
backtrack[4][14] <= nxt_backtrack[4][14];
backtrack[4][15] <= nxt_backtrack[4][15];
backtrack[4][16] <= nxt_backtrack[4][16];
backtrack[4][17] <= nxt_backtrack[4][17];
backtrack[4][18] <= nxt_backtrack[4][18];
backtrack[4][19] <= nxt_backtrack[4][19];
backtrack[5][0] <= nxt_backtrack[5][0];
backtrack[5][1] <= nxt_backtrack[5][1];
backtrack[5][2] <= nxt_backtrack[5][2];
backtrack[5][3] <= nxt_backtrack[5][3];
backtrack[5][4] <= nxt_backtrack[5][4];
backtrack[5][5] <= nxt_backtrack[5][5];
backtrack[5][6] <= nxt_backtrack[5][6];
backtrack[5][7] <= nxt_backtrack[5][7];
backtrack[5][8] <= nxt_backtrack[5][8];
backtrack[5][9] <= nxt_backtrack[5][9];
backtrack[5][10] <= nxt_backtrack[5][10];
backtrack[5][11] <= nxt_backtrack[5][11];
backtrack[5][12] <= nxt_backtrack[5][12];
backtrack[5][13] <= nxt_backtrack[5][13];
backtrack[5][14] <= nxt_backtrack[5][14];
backtrack[5][15] <= nxt_backtrack[5][15];
backtrack[5][16] <= nxt_backtrack[5][16];
backtrack[5][17] <= nxt_backtrack[5][17];
backtrack[5][18] <= nxt_backtrack[5][18];
backtrack[5][19] <= nxt_backtrack[5][19];
backtrack[6][0] <= nxt_backtrack[6][0];
backtrack[6][1] <= nxt_backtrack[6][1];
backtrack[6][2] <= nxt_backtrack[6][2];
backtrack[6][3] <= nxt_backtrack[6][3];
backtrack[6][4] <= nxt_backtrack[6][4];
backtrack[6][5] <= nxt_backtrack[6][5];
backtrack[6][6] <= nxt_backtrack[6][6];
backtrack[6][7] <= nxt_backtrack[6][7];
backtrack[6][8] <= nxt_backtrack[6][8];
backtrack[6][9] <= nxt_backtrack[6][9];
backtrack[6][10] <= nxt_backtrack[6][10];
backtrack[6][11] <= nxt_backtrack[6][11];
backtrack[6][12] <= nxt_backtrack[6][12];
backtrack[6][13] <= nxt_backtrack[6][13];
backtrack[6][14] <= nxt_backtrack[6][14];
backtrack[6][15] <= nxt_backtrack[6][15];
backtrack[6][16] <= nxt_backtrack[6][16];
backtrack[6][17] <= nxt_backtrack[6][17];
backtrack[6][18] <= nxt_backtrack[6][18];
backtrack[6][19] <= nxt_backtrack[6][19];
backtrack[7][0] <= nxt_backtrack[7][0];
backtrack[7][1] <= nxt_backtrack[7][1];
backtrack[7][2] <= nxt_backtrack[7][2];
backtrack[7][3] <= nxt_backtrack[7][3];
backtrack[7][4] <= nxt_backtrack[7][4];
backtrack[7][5] <= nxt_backtrack[7][5];
backtrack[7][6] <= nxt_backtrack[7][6];
backtrack[7][7] <= nxt_backtrack[7][7];
backtrack[7][8] <= nxt_backtrack[7][8];
backtrack[7][9] <= nxt_backtrack[7][9];
backtrack[7][10] <= nxt_backtrack[7][10];
backtrack[7][11] <= nxt_backtrack[7][11];
backtrack[7][12] <= nxt_backtrack[7][12];
backtrack[7][13] <= nxt_backtrack[7][13];
backtrack[7][14] <= nxt_backtrack[7][14];
backtrack[7][15] <= nxt_backtrack[7][15];
backtrack[7][16] <= nxt_backtrack[7][16];
backtrack[7][17] <= nxt_backtrack[7][17];
backtrack[7][18] <= nxt_backtrack[7][18];
backtrack[7][19] <= nxt_backtrack[7][19];
backtrack[8][0] <= nxt_backtrack[8][0];
backtrack[8][1] <= nxt_backtrack[8][1];
backtrack[8][2] <= nxt_backtrack[8][2];
backtrack[8][3] <= nxt_backtrack[8][3];
backtrack[8][4] <= nxt_backtrack[8][4];
backtrack[8][5] <= nxt_backtrack[8][5];
backtrack[8][6] <= nxt_backtrack[8][6];
backtrack[8][7] <= nxt_backtrack[8][7];
backtrack[8][8] <= nxt_backtrack[8][8];
backtrack[8][9] <= nxt_backtrack[8][9];
backtrack[8][10] <= nxt_backtrack[8][10];
backtrack[8][11] <= nxt_backtrack[8][11];
backtrack[8][12] <= nxt_backtrack[8][12];
backtrack[8][13] <= nxt_backtrack[8][13];
backtrack[8][14] <= nxt_backtrack[8][14];
backtrack[8][15] <= nxt_backtrack[8][15];
backtrack[8][16] <= nxt_backtrack[8][16];
backtrack[8][17] <= nxt_backtrack[8][17];
backtrack[8][18] <= nxt_backtrack[8][18];
backtrack[8][19] <= nxt_backtrack[8][19];
backtrack[9][0] <= nxt_backtrack[9][0];
backtrack[9][1] <= nxt_backtrack[9][1];
backtrack[9][2] <= nxt_backtrack[9][2];
backtrack[9][3] <= nxt_backtrack[9][3];
backtrack[9][4] <= nxt_backtrack[9][4];
backtrack[9][5] <= nxt_backtrack[9][5];
backtrack[9][6] <= nxt_backtrack[9][6];
backtrack[9][7] <= nxt_backtrack[9][7];
backtrack[9][8] <= nxt_backtrack[9][8];
backtrack[9][9] <= nxt_backtrack[9][9];
backtrack[9][10] <= nxt_backtrack[9][10];
backtrack[9][11] <= nxt_backtrack[9][11];
backtrack[9][12] <= nxt_backtrack[9][12];
backtrack[9][13] <= nxt_backtrack[9][13];
backtrack[9][14] <= nxt_backtrack[9][14];
backtrack[9][15] <= nxt_backtrack[9][15];
backtrack[9][16] <= nxt_backtrack[9][16];
backtrack[9][17] <= nxt_backtrack[9][17];
backtrack[9][18] <= nxt_backtrack[9][18];
backtrack[9][19] <= nxt_backtrack[9][19];
end
endtask
task shift_shortest_dist;
begin
shortest_dist[0][0] <= nxt_shortest_dist[0][0];
shortest_dist[0][1] <= nxt_shortest_dist[0][1];
shortest_dist[0][2] <= nxt_shortest_dist[0][2];
shortest_dist[0][3] <= nxt_shortest_dist[0][3];
shortest_dist[0][4] <= nxt_shortest_dist[0][4];
shortest_dist[0][5] <= nxt_shortest_dist[0][5];
shortest_dist[0][6] <= nxt_shortest_dist[0][6];
shortest_dist[0][7] <= nxt_shortest_dist[0][7];
shortest_dist[0][8] <= nxt_shortest_dist[0][8];
shortest_dist[0][9] <= nxt_shortest_dist[0][9];
shortest_dist[0][10] <= nxt_shortest_dist[0][10];
shortest_dist[0][11] <= nxt_shortest_dist[0][11];
shortest_dist[0][12] <= nxt_shortest_dist[0][12];
shortest_dist[0][13] <= nxt_shortest_dist[0][13];
shortest_dist[0][14] <= nxt_shortest_dist[0][14];
shortest_dist[0][15] <= nxt_shortest_dist[0][15];
shortest_dist[0][16] <= nxt_shortest_dist[0][16];
shortest_dist[0][17] <= nxt_shortest_dist[0][17];
shortest_dist[0][18] <= nxt_shortest_dist[0][18];
shortest_dist[0][19] <= nxt_shortest_dist[0][19];
shortest_dist[1][0] <= nxt_shortest_dist[1][0];
shortest_dist[1][1] <= nxt_shortest_dist[1][1];
shortest_dist[1][2] <= nxt_shortest_dist[1][2];
shortest_dist[1][3] <= nxt_shortest_dist[1][3];
shortest_dist[1][4] <= nxt_shortest_dist[1][4];
shortest_dist[1][5] <= nxt_shortest_dist[1][5];
shortest_dist[1][6] <= nxt_shortest_dist[1][6];
shortest_dist[1][7] <= nxt_shortest_dist[1][7];
shortest_dist[1][8] <= nxt_shortest_dist[1][8];
shortest_dist[1][9] <= nxt_shortest_dist[1][9];
shortest_dist[1][10] <= nxt_shortest_dist[1][10];
shortest_dist[1][11] <= nxt_shortest_dist[1][11];
shortest_dist[1][12] <= nxt_shortest_dist[1][12];
shortest_dist[1][13] <= nxt_shortest_dist[1][13];
shortest_dist[1][14] <= nxt_shortest_dist[1][14];
shortest_dist[1][15] <= nxt_shortest_dist[1][15];
shortest_dist[1][16] <= nxt_shortest_dist[1][16];
shortest_dist[1][17] <= nxt_shortest_dist[1][17];
shortest_dist[1][18] <= nxt_shortest_dist[1][18];
shortest_dist[1][19] <= nxt_shortest_dist[1][19];
shortest_dist[2][0] <= nxt_shortest_dist[2][0];
shortest_dist[2][1] <= nxt_shortest_dist[2][1];
shortest_dist[2][2] <= nxt_shortest_dist[2][2];
shortest_dist[2][3] <= nxt_shortest_dist[2][3];
shortest_dist[2][4] <= nxt_shortest_dist[2][4];
shortest_dist[2][5] <= nxt_shortest_dist[2][5];
shortest_dist[2][6] <= nxt_shortest_dist[2][6];
shortest_dist[2][7] <= nxt_shortest_dist[2][7];
shortest_dist[2][8] <= nxt_shortest_dist[2][8];
shortest_dist[2][9] <= nxt_shortest_dist[2][9];
shortest_dist[2][10] <= nxt_shortest_dist[2][10];
shortest_dist[2][11] <= nxt_shortest_dist[2][11];
shortest_dist[2][12] <= nxt_shortest_dist[2][12];
shortest_dist[2][13] <= nxt_shortest_dist[2][13];
shortest_dist[2][14] <= nxt_shortest_dist[2][14];
shortest_dist[2][15] <= nxt_shortest_dist[2][15];
shortest_dist[2][16] <= nxt_shortest_dist[2][16];
shortest_dist[2][17] <= nxt_shortest_dist[2][17];
shortest_dist[2][18] <= nxt_shortest_dist[2][18];
shortest_dist[2][19] <= nxt_shortest_dist[2][19];
shortest_dist[3][0] <= nxt_shortest_dist[3][0];
shortest_dist[3][1] <= nxt_shortest_dist[3][1];
shortest_dist[3][2] <= nxt_shortest_dist[3][2];
shortest_dist[3][3] <= nxt_shortest_dist[3][3];
shortest_dist[3][4] <= nxt_shortest_dist[3][4];
shortest_dist[3][5] <= nxt_shortest_dist[3][5];
shortest_dist[3][6] <= nxt_shortest_dist[3][6];
shortest_dist[3][7] <= nxt_shortest_dist[3][7];
shortest_dist[3][8] <= nxt_shortest_dist[3][8];
shortest_dist[3][9] <= nxt_shortest_dist[3][9];
shortest_dist[3][10] <= nxt_shortest_dist[3][10];
shortest_dist[3][11] <= nxt_shortest_dist[3][11];
shortest_dist[3][12] <= nxt_shortest_dist[3][12];
shortest_dist[3][13] <= nxt_shortest_dist[3][13];
shortest_dist[3][14] <= nxt_shortest_dist[3][14];
shortest_dist[3][15] <= nxt_shortest_dist[3][15];
shortest_dist[3][16] <= nxt_shortest_dist[3][16];
shortest_dist[3][17] <= nxt_shortest_dist[3][17];
shortest_dist[3][18] <= nxt_shortest_dist[3][18];
shortest_dist[3][19] <= nxt_shortest_dist[3][19];
shortest_dist[4][0] <= nxt_shortest_dist[4][0];
shortest_dist[4][1] <= nxt_shortest_dist[4][1];
shortest_dist[4][2] <= nxt_shortest_dist[4][2];
shortest_dist[4][3] <= nxt_shortest_dist[4][3];
shortest_dist[4][4] <= nxt_shortest_dist[4][4];
shortest_dist[4][5] <= nxt_shortest_dist[4][5];
shortest_dist[4][6] <= nxt_shortest_dist[4][6];
shortest_dist[4][7] <= nxt_shortest_dist[4][7];
shortest_dist[4][8] <= nxt_shortest_dist[4][8];
shortest_dist[4][9] <= nxt_shortest_dist[4][9];
shortest_dist[4][10] <= nxt_shortest_dist[4][10];
shortest_dist[4][11] <= nxt_shortest_dist[4][11];
shortest_dist[4][12] <= nxt_shortest_dist[4][12];
shortest_dist[4][13] <= nxt_shortest_dist[4][13];
shortest_dist[4][14] <= nxt_shortest_dist[4][14];
shortest_dist[4][15] <= nxt_shortest_dist[4][15];
shortest_dist[4][16] <= nxt_shortest_dist[4][16];
shortest_dist[4][17] <= nxt_shortest_dist[4][17];
shortest_dist[4][18] <= nxt_shortest_dist[4][18];
shortest_dist[4][19] <= nxt_shortest_dist[4][19];
shortest_dist[5][0] <= nxt_shortest_dist[5][0];
shortest_dist[5][1] <= nxt_shortest_dist[5][1];
shortest_dist[5][2] <= nxt_shortest_dist[5][2];
shortest_dist[5][3] <= nxt_shortest_dist[5][3];
shortest_dist[5][4] <= nxt_shortest_dist[5][4];
shortest_dist[5][5] <= nxt_shortest_dist[5][5];
shortest_dist[5][6] <= nxt_shortest_dist[5][6];
shortest_dist[5][7] <= nxt_shortest_dist[5][7];
shortest_dist[5][8] <= nxt_shortest_dist[5][8];
shortest_dist[5][9] <= nxt_shortest_dist[5][9];
shortest_dist[5][10] <= nxt_shortest_dist[5][10];
shortest_dist[5][11] <= nxt_shortest_dist[5][11];
shortest_dist[5][12] <= nxt_shortest_dist[5][12];
shortest_dist[5][13] <= nxt_shortest_dist[5][13];
shortest_dist[5][14] <= nxt_shortest_dist[5][14];
shortest_dist[5][15] <= nxt_shortest_dist[5][15];
shortest_dist[5][16] <= nxt_shortest_dist[5][16];
shortest_dist[5][17] <= nxt_shortest_dist[5][17];
shortest_dist[5][18] <= nxt_shortest_dist[5][18];
shortest_dist[5][19] <= nxt_shortest_dist[5][19];
shortest_dist[6][0] <= nxt_shortest_dist[6][0];
shortest_dist[6][1] <= nxt_shortest_dist[6][1];
shortest_dist[6][2] <= nxt_shortest_dist[6][2];
shortest_dist[6][3] <= nxt_shortest_dist[6][3];
shortest_dist[6][4] <= nxt_shortest_dist[6][4];
shortest_dist[6][5] <= nxt_shortest_dist[6][5];
shortest_dist[6][6] <= nxt_shortest_dist[6][6];
shortest_dist[6][7] <= nxt_shortest_dist[6][7];
shortest_dist[6][8] <= nxt_shortest_dist[6][8];
shortest_dist[6][9] <= nxt_shortest_dist[6][9];
shortest_dist[6][10] <= nxt_shortest_dist[6][10];
shortest_dist[6][11] <= nxt_shortest_dist[6][11];
shortest_dist[6][12] <= nxt_shortest_dist[6][12];
shortest_dist[6][13] <= nxt_shortest_dist[6][13];
shortest_dist[6][14] <= nxt_shortest_dist[6][14];
shortest_dist[6][15] <= nxt_shortest_dist[6][15];
shortest_dist[6][16] <= nxt_shortest_dist[6][16];
shortest_dist[6][17] <= nxt_shortest_dist[6][17];
shortest_dist[6][18] <= nxt_shortest_dist[6][18];
shortest_dist[6][19] <= nxt_shortest_dist[6][19];
shortest_dist[7][0] <= nxt_shortest_dist[7][0];
shortest_dist[7][1] <= nxt_shortest_dist[7][1];
shortest_dist[7][2] <= nxt_shortest_dist[7][2];
shortest_dist[7][3] <= nxt_shortest_dist[7][3];
shortest_dist[7][4] <= nxt_shortest_dist[7][4];
shortest_dist[7][5] <= nxt_shortest_dist[7][5];
shortest_dist[7][6] <= nxt_shortest_dist[7][6];
shortest_dist[7][7] <= nxt_shortest_dist[7][7];
shortest_dist[7][8] <= nxt_shortest_dist[7][8];
shortest_dist[7][9] <= nxt_shortest_dist[7][9];
shortest_dist[7][10] <= nxt_shortest_dist[7][10];
shortest_dist[7][11] <= nxt_shortest_dist[7][11];
shortest_dist[7][12] <= nxt_shortest_dist[7][12];
shortest_dist[7][13] <= nxt_shortest_dist[7][13];
shortest_dist[7][14] <= nxt_shortest_dist[7][14];
shortest_dist[7][15] <= nxt_shortest_dist[7][15];
shortest_dist[7][16] <= nxt_shortest_dist[7][16];
shortest_dist[7][17] <= nxt_shortest_dist[7][17];
shortest_dist[7][18] <= nxt_shortest_dist[7][18];
shortest_dist[7][19] <= nxt_shortest_dist[7][19];
shortest_dist[8][0] <= nxt_shortest_dist[8][0];
shortest_dist[8][1] <= nxt_shortest_dist[8][1];
shortest_dist[8][2] <= nxt_shortest_dist[8][2];
shortest_dist[8][3] <= nxt_shortest_dist[8][3];
shortest_dist[8][4] <= nxt_shortest_dist[8][4];
shortest_dist[8][5] <= nxt_shortest_dist[8][5];
shortest_dist[8][6] <= nxt_shortest_dist[8][6];
shortest_dist[8][7] <= nxt_shortest_dist[8][7];
shortest_dist[8][8] <= nxt_shortest_dist[8][8];
shortest_dist[8][9] <= nxt_shortest_dist[8][9];
shortest_dist[8][10] <= nxt_shortest_dist[8][10];
shortest_dist[8][11] <= nxt_shortest_dist[8][11];
shortest_dist[8][12] <= nxt_shortest_dist[8][12];
shortest_dist[8][13] <= nxt_shortest_dist[8][13];
shortest_dist[8][14] <= nxt_shortest_dist[8][14];
shortest_dist[8][15] <= nxt_shortest_dist[8][15];
shortest_dist[8][16] <= nxt_shortest_dist[8][16];
shortest_dist[8][17] <= nxt_shortest_dist[8][17];
shortest_dist[8][18] <= nxt_shortest_dist[8][18];
shortest_dist[8][19] <= nxt_shortest_dist[8][19];
shortest_dist[9][0] <= nxt_shortest_dist[9][0];
shortest_dist[9][1] <= nxt_shortest_dist[9][1];
shortest_dist[9][2] <= nxt_shortest_dist[9][2];
shortest_dist[9][3] <= nxt_shortest_dist[9][3];
shortest_dist[9][4] <= nxt_shortest_dist[9][4];
shortest_dist[9][5] <= nxt_shortest_dist[9][5];
shortest_dist[9][6] <= nxt_shortest_dist[9][6];
shortest_dist[9][7] <= nxt_shortest_dist[9][7];
shortest_dist[9][8] <= nxt_shortest_dist[9][8];
shortest_dist[9][9] <= nxt_shortest_dist[9][9];
shortest_dist[9][10] <= nxt_shortest_dist[9][10];
shortest_dist[9][11] <= nxt_shortest_dist[9][11];
shortest_dist[9][12] <= nxt_shortest_dist[9][12];
shortest_dist[9][13] <= nxt_shortest_dist[9][13];
shortest_dist[9][14] <= nxt_shortest_dist[9][14];
shortest_dist[9][15] <= nxt_shortest_dist[9][15];
shortest_dist[9][16] <= nxt_shortest_dist[9][16];
shortest_dist[9][17] <= nxt_shortest_dist[9][17];
shortest_dist[9][18] <= nxt_shortest_dist[9][18];
shortest_dist[9][19] <= nxt_shortest_dist[9][19];
end
endtask
task shift_nxt_backtrack;
begin
nxt_backtrack[0][0] <= backtrack[0][0];
nxt_backtrack[0][1] <= backtrack[0][1];
nxt_backtrack[0][2] <= backtrack[0][2];
nxt_backtrack[0][3] <= backtrack[0][3];
nxt_backtrack[0][4] <= backtrack[0][4];
nxt_backtrack[0][5] <= backtrack[0][5];
nxt_backtrack[0][6] <= backtrack[0][6];
nxt_backtrack[0][7] <= backtrack[0][7];
nxt_backtrack[0][8] <= backtrack[0][8];
nxt_backtrack[0][9] <= backtrack[0][9];
nxt_backtrack[0][10] <= backtrack[0][10];
nxt_backtrack[0][11] <= backtrack[0][11];
nxt_backtrack[0][12] <= backtrack[0][12];
nxt_backtrack[0][13] <= backtrack[0][13];
nxt_backtrack[0][14] <= backtrack[0][14];
nxt_backtrack[0][15] <= backtrack[0][15];
nxt_backtrack[0][16] <= backtrack[0][16];
nxt_backtrack[0][17] <= backtrack[0][17];
nxt_backtrack[0][18] <= backtrack[0][18];
nxt_backtrack[0][19] <= backtrack[0][19];
nxt_backtrack[1][0] <= backtrack[1][0];
nxt_backtrack[1][1] <= backtrack[1][1];
nxt_backtrack[1][2] <= backtrack[1][2];
nxt_backtrack[1][3] <= backtrack[1][3];
nxt_backtrack[1][4] <= backtrack[1][4];
nxt_backtrack[1][5] <= backtrack[1][5];
nxt_backtrack[1][6] <= backtrack[1][6];
nxt_backtrack[1][7] <= backtrack[1][7];
nxt_backtrack[1][8] <= backtrack[1][8];
nxt_backtrack[1][9] <= backtrack[1][9];
nxt_backtrack[1][10] <= backtrack[1][10];
nxt_backtrack[1][11] <= backtrack[1][11];
nxt_backtrack[1][12] <= backtrack[1][12];
nxt_backtrack[1][13] <= backtrack[1][13];
nxt_backtrack[1][14] <= backtrack[1][14];
nxt_backtrack[1][15] <= backtrack[1][15];
nxt_backtrack[1][16] <= backtrack[1][16];
nxt_backtrack[1][17] <= backtrack[1][17];
nxt_backtrack[1][18] <= backtrack[1][18];
nxt_backtrack[1][19] <= backtrack[1][19];
nxt_backtrack[2][0] <= backtrack[2][0];
nxt_backtrack[2][1] <= backtrack[2][1];
nxt_backtrack[2][2] <= backtrack[2][2];
nxt_backtrack[2][3] <= backtrack[2][3];
nxt_backtrack[2][4] <= backtrack[2][4];
nxt_backtrack[2][5] <= backtrack[2][5];
nxt_backtrack[2][6] <= backtrack[2][6];
nxt_backtrack[2][7] <= backtrack[2][7];
nxt_backtrack[2][8] <= backtrack[2][8];
nxt_backtrack[2][9] <= backtrack[2][9];
nxt_backtrack[2][10] <= backtrack[2][10];
nxt_backtrack[2][11] <= backtrack[2][11];
nxt_backtrack[2][12] <= backtrack[2][12];
nxt_backtrack[2][13] <= backtrack[2][13];
nxt_backtrack[2][14] <= backtrack[2][14];
nxt_backtrack[2][15] <= backtrack[2][15];
nxt_backtrack[2][16] <= backtrack[2][16];
nxt_backtrack[2][17] <= backtrack[2][17];
nxt_backtrack[2][18] <= backtrack[2][18];
nxt_backtrack[2][19] <= backtrack[2][19];
nxt_backtrack[3][0] <= backtrack[3][0];
nxt_backtrack[3][1] <= backtrack[3][1];
nxt_backtrack[3][2] <= backtrack[3][2];
nxt_backtrack[3][3] <= backtrack[3][3];
nxt_backtrack[3][4] <= backtrack[3][4];
nxt_backtrack[3][5] <= backtrack[3][5];
nxt_backtrack[3][6] <= backtrack[3][6];
nxt_backtrack[3][7] <= backtrack[3][7];
nxt_backtrack[3][8] <= backtrack[3][8];
nxt_backtrack[3][9] <= backtrack[3][9];
nxt_backtrack[3][10] <= backtrack[3][10];
nxt_backtrack[3][11] <= backtrack[3][11];
nxt_backtrack[3][12] <= backtrack[3][12];
nxt_backtrack[3][13] <= backtrack[3][13];
nxt_backtrack[3][14] <= backtrack[3][14];
nxt_backtrack[3][15] <= backtrack[3][15];
nxt_backtrack[3][16] <= backtrack[3][16];
nxt_backtrack[3][17] <= backtrack[3][17];
nxt_backtrack[3][18] <= backtrack[3][18];
nxt_backtrack[3][19] <= backtrack[3][19];
nxt_backtrack[4][0] <= backtrack[4][0];
nxt_backtrack[4][1] <= backtrack[4][1];
nxt_backtrack[4][2] <= backtrack[4][2];
nxt_backtrack[4][3] <= backtrack[4][3];
nxt_backtrack[4][4] <= backtrack[4][4];
nxt_backtrack[4][5] <= backtrack[4][5];
nxt_backtrack[4][6] <= backtrack[4][6];
nxt_backtrack[4][7] <= backtrack[4][7];
nxt_backtrack[4][8] <= backtrack[4][8];
nxt_backtrack[4][9] <= backtrack[4][9];
nxt_backtrack[4][10] <= backtrack[4][10];
nxt_backtrack[4][11] <= backtrack[4][11];
nxt_backtrack[4][12] <= backtrack[4][12];
nxt_backtrack[4][13] <= backtrack[4][13];
nxt_backtrack[4][14] <= backtrack[4][14];
nxt_backtrack[4][15] <= backtrack[4][15];
nxt_backtrack[4][16] <= backtrack[4][16];
nxt_backtrack[4][17] <= backtrack[4][17];
nxt_backtrack[4][18] <= backtrack[4][18];
nxt_backtrack[4][19] <= backtrack[4][19];
nxt_backtrack[5][0] <= backtrack[5][0];
nxt_backtrack[5][1] <= backtrack[5][1];
nxt_backtrack[5][2] <= backtrack[5][2];
nxt_backtrack[5][3] <= backtrack[5][3];
nxt_backtrack[5][4] <= backtrack[5][4];
nxt_backtrack[5][5] <= backtrack[5][5];
nxt_backtrack[5][6] <= backtrack[5][6];
nxt_backtrack[5][7] <= backtrack[5][7];
nxt_backtrack[5][8] <= backtrack[5][8];
nxt_backtrack[5][9] <= backtrack[5][9];
nxt_backtrack[5][10] <= backtrack[5][10];
nxt_backtrack[5][11] <= backtrack[5][11];
nxt_backtrack[5][12] <= backtrack[5][12];
nxt_backtrack[5][13] <= backtrack[5][13];
nxt_backtrack[5][14] <= backtrack[5][14];
nxt_backtrack[5][15] <= backtrack[5][15];
nxt_backtrack[5][16] <= backtrack[5][16];
nxt_backtrack[5][17] <= backtrack[5][17];
nxt_backtrack[5][18] <= backtrack[5][18];
nxt_backtrack[5][19] <= backtrack[5][19];
nxt_backtrack[6][0] <= backtrack[6][0];
nxt_backtrack[6][1] <= backtrack[6][1];
nxt_backtrack[6][2] <= backtrack[6][2];
nxt_backtrack[6][3] <= backtrack[6][3];
nxt_backtrack[6][4] <= backtrack[6][4];
nxt_backtrack[6][5] <= backtrack[6][5];
nxt_backtrack[6][6] <= backtrack[6][6];
nxt_backtrack[6][7] <= backtrack[6][7];
nxt_backtrack[6][8] <= backtrack[6][8];
nxt_backtrack[6][9] <= backtrack[6][9];
nxt_backtrack[6][10] <= backtrack[6][10];
nxt_backtrack[6][11] <= backtrack[6][11];
nxt_backtrack[6][12] <= backtrack[6][12];
nxt_backtrack[6][13] <= backtrack[6][13];
nxt_backtrack[6][14] <= backtrack[6][14];
nxt_backtrack[6][15] <= backtrack[6][15];
nxt_backtrack[6][16] <= backtrack[6][16];
nxt_backtrack[6][17] <= backtrack[6][17];
nxt_backtrack[6][18] <= backtrack[6][18];
nxt_backtrack[6][19] <= backtrack[6][19];
nxt_backtrack[7][0] <= backtrack[7][0];
nxt_backtrack[7][1] <= backtrack[7][1];
nxt_backtrack[7][2] <= backtrack[7][2];
nxt_backtrack[7][3] <= backtrack[7][3];
nxt_backtrack[7][4] <= backtrack[7][4];
nxt_backtrack[7][5] <= backtrack[7][5];
nxt_backtrack[7][6] <= backtrack[7][6];
nxt_backtrack[7][7] <= backtrack[7][7];
nxt_backtrack[7][8] <= backtrack[7][8];
nxt_backtrack[7][9] <= backtrack[7][9];
nxt_backtrack[7][10] <= backtrack[7][10];
nxt_backtrack[7][11] <= backtrack[7][11];
nxt_backtrack[7][12] <= backtrack[7][12];
nxt_backtrack[7][13] <= backtrack[7][13];
nxt_backtrack[7][14] <= backtrack[7][14];
nxt_backtrack[7][15] <= backtrack[7][15];
nxt_backtrack[7][16] <= backtrack[7][16];
nxt_backtrack[7][17] <= backtrack[7][17];
nxt_backtrack[7][18] <= backtrack[7][18];
nxt_backtrack[7][19] <= backtrack[7][19];
nxt_backtrack[8][0] <= backtrack[8][0];
nxt_backtrack[8][1] <= backtrack[8][1];
nxt_backtrack[8][2] <= backtrack[8][2];
nxt_backtrack[8][3] <= backtrack[8][3];
nxt_backtrack[8][4] <= backtrack[8][4];
nxt_backtrack[8][5] <= backtrack[8][5];
nxt_backtrack[8][6] <= backtrack[8][6];
nxt_backtrack[8][7] <= backtrack[8][7];
nxt_backtrack[8][8] <= backtrack[8][8];
nxt_backtrack[8][9] <= backtrack[8][9];
nxt_backtrack[8][10] <= backtrack[8][10];
nxt_backtrack[8][11] <= backtrack[8][11];
nxt_backtrack[8][12] <= backtrack[8][12];
nxt_backtrack[8][13] <= backtrack[8][13];
nxt_backtrack[8][14] <= backtrack[8][14];
nxt_backtrack[8][15] <= backtrack[8][15];
nxt_backtrack[8][16] <= backtrack[8][16];
nxt_backtrack[8][17] <= backtrack[8][17];
nxt_backtrack[8][18] <= backtrack[8][18];
nxt_backtrack[8][19] <= backtrack[8][19];
nxt_backtrack[9][0] <= backtrack[9][0];
nxt_backtrack[9][1] <= backtrack[9][1];
nxt_backtrack[9][2] <= backtrack[9][2];
nxt_backtrack[9][3] <= backtrack[9][3];
nxt_backtrack[9][4] <= backtrack[9][4];
nxt_backtrack[9][5] <= backtrack[9][5];
nxt_backtrack[9][6] <= backtrack[9][6];
nxt_backtrack[9][7] <= backtrack[9][7];
nxt_backtrack[9][8] <= backtrack[9][8];
nxt_backtrack[9][9] <= backtrack[9][9];
nxt_backtrack[9][10] <= backtrack[9][10];
nxt_backtrack[9][11] <= backtrack[9][11];
nxt_backtrack[9][12] <= backtrack[9][12];
nxt_backtrack[9][13] <= backtrack[9][13];
nxt_backtrack[9][14] <= backtrack[9][14];
nxt_backtrack[9][15] <= backtrack[9][15];
nxt_backtrack[9][16] <= backtrack[9][16];
nxt_backtrack[9][17] <= backtrack[9][17];
nxt_backtrack[9][18] <= backtrack[9][18];
nxt_backtrack[9][19] <= backtrack[9][19];
end
endtask
task shift_nxt_shortest_dist;
begin
nxt_shortest_dist[0][0] <= shortest_dist[0][0];
nxt_shortest_dist[0][1] <= shortest_dist[0][1];
nxt_shortest_dist[0][2] <= shortest_dist[0][2];
nxt_shortest_dist[0][3] <= shortest_dist[0][3];
nxt_shortest_dist[0][4] <= shortest_dist[0][4];
nxt_shortest_dist[0][5] <= shortest_dist[0][5];
nxt_shortest_dist[0][6] <= shortest_dist[0][6];
nxt_shortest_dist[0][7] <= shortest_dist[0][7];
nxt_shortest_dist[0][8] <= shortest_dist[0][8];
nxt_shortest_dist[0][9] <= shortest_dist[0][9];
nxt_shortest_dist[0][10] <= shortest_dist[0][10];
nxt_shortest_dist[0][11] <= shortest_dist[0][11];
nxt_shortest_dist[0][12] <= shortest_dist[0][12];
nxt_shortest_dist[0][13] <= shortest_dist[0][13];
nxt_shortest_dist[0][14] <= shortest_dist[0][14];
nxt_shortest_dist[0][15] <= shortest_dist[0][15];
nxt_shortest_dist[0][16] <= shortest_dist[0][16];
nxt_shortest_dist[0][17] <= shortest_dist[0][17];
nxt_shortest_dist[0][18] <= shortest_dist[0][18];
nxt_shortest_dist[0][19] <= shortest_dist[0][19];
nxt_shortest_dist[1][0] <= shortest_dist[1][0];
nxt_shortest_dist[1][1] <= shortest_dist[1][1];
nxt_shortest_dist[1][2] <= shortest_dist[1][2];
nxt_shortest_dist[1][3] <= shortest_dist[1][3];
nxt_shortest_dist[1][4] <= shortest_dist[1][4];
nxt_shortest_dist[1][5] <= shortest_dist[1][5];
nxt_shortest_dist[1][6] <= shortest_dist[1][6];
nxt_shortest_dist[1][7] <= shortest_dist[1][7];
nxt_shortest_dist[1][8] <= shortest_dist[1][8];
nxt_shortest_dist[1][9] <= shortest_dist[1][9];
nxt_shortest_dist[1][10] <= shortest_dist[1][10];
nxt_shortest_dist[1][11] <= shortest_dist[1][11];
nxt_shortest_dist[1][12] <= shortest_dist[1][12];
nxt_shortest_dist[1][13] <= shortest_dist[1][13];
nxt_shortest_dist[1][14] <= shortest_dist[1][14];
nxt_shortest_dist[1][15] <= shortest_dist[1][15];
nxt_shortest_dist[1][16] <= shortest_dist[1][16];
nxt_shortest_dist[1][17] <= shortest_dist[1][17];
nxt_shortest_dist[1][18] <= shortest_dist[1][18];
nxt_shortest_dist[1][19] <= shortest_dist[1][19];
nxt_shortest_dist[2][0] <= shortest_dist[2][0];
nxt_shortest_dist[2][1] <= shortest_dist[2][1];
nxt_shortest_dist[2][2] <= shortest_dist[2][2];
nxt_shortest_dist[2][3] <= shortest_dist[2][3];
nxt_shortest_dist[2][4] <= shortest_dist[2][4];
nxt_shortest_dist[2][5] <= shortest_dist[2][5];
nxt_shortest_dist[2][6] <= shortest_dist[2][6];
nxt_shortest_dist[2][7] <= shortest_dist[2][7];
nxt_shortest_dist[2][8] <= shortest_dist[2][8];
nxt_shortest_dist[2][9] <= shortest_dist[2][9];
nxt_shortest_dist[2][10] <= shortest_dist[2][10];
nxt_shortest_dist[2][11] <= shortest_dist[2][11];
nxt_shortest_dist[2][12] <= shortest_dist[2][12];
nxt_shortest_dist[2][13] <= shortest_dist[2][13];
nxt_shortest_dist[2][14] <= shortest_dist[2][14];
nxt_shortest_dist[2][15] <= shortest_dist[2][15];
nxt_shortest_dist[2][16] <= shortest_dist[2][16];
nxt_shortest_dist[2][17] <= shortest_dist[2][17];
nxt_shortest_dist[2][18] <= shortest_dist[2][18];
nxt_shortest_dist[2][19] <= shortest_dist[2][19];
nxt_shortest_dist[3][0] <= shortest_dist[3][0];
nxt_shortest_dist[3][1] <= shortest_dist[3][1];
nxt_shortest_dist[3][2] <= shortest_dist[3][2];
nxt_shortest_dist[3][3] <= shortest_dist[3][3];
nxt_shortest_dist[3][4] <= shortest_dist[3][4];
nxt_shortest_dist[3][5] <= shortest_dist[3][5];
nxt_shortest_dist[3][6] <= shortest_dist[3][6];
nxt_shortest_dist[3][7] <= shortest_dist[3][7];
nxt_shortest_dist[3][8] <= shortest_dist[3][8];
nxt_shortest_dist[3][9] <= shortest_dist[3][9];
nxt_shortest_dist[3][10] <= shortest_dist[3][10];
nxt_shortest_dist[3][11] <= shortest_dist[3][11];
nxt_shortest_dist[3][12] <= shortest_dist[3][12];
nxt_shortest_dist[3][13] <= shortest_dist[3][13];
nxt_shortest_dist[3][14] <= shortest_dist[3][14];
nxt_shortest_dist[3][15] <= shortest_dist[3][15];
nxt_shortest_dist[3][16] <= shortest_dist[3][16];
nxt_shortest_dist[3][17] <= shortest_dist[3][17];
nxt_shortest_dist[3][18] <= shortest_dist[3][18];
nxt_shortest_dist[3][19] <= shortest_dist[3][19];
nxt_shortest_dist[4][0] <= shortest_dist[4][0];
nxt_shortest_dist[4][1] <= shortest_dist[4][1];
nxt_shortest_dist[4][2] <= shortest_dist[4][2];
nxt_shortest_dist[4][3] <= shortest_dist[4][3];
nxt_shortest_dist[4][4] <= shortest_dist[4][4];
nxt_shortest_dist[4][5] <= shortest_dist[4][5];
nxt_shortest_dist[4][6] <= shortest_dist[4][6];
nxt_shortest_dist[4][7] <= shortest_dist[4][7];
nxt_shortest_dist[4][8] <= shortest_dist[4][8];
nxt_shortest_dist[4][9] <= shortest_dist[4][9];
nxt_shortest_dist[4][10] <= shortest_dist[4][10];
nxt_shortest_dist[4][11] <= shortest_dist[4][11];
nxt_shortest_dist[4][12] <= shortest_dist[4][12];
nxt_shortest_dist[4][13] <= shortest_dist[4][13];
nxt_shortest_dist[4][14] <= shortest_dist[4][14];
nxt_shortest_dist[4][15] <= shortest_dist[4][15];
nxt_shortest_dist[4][16] <= shortest_dist[4][16];
nxt_shortest_dist[4][17] <= shortest_dist[4][17];
nxt_shortest_dist[4][18] <= shortest_dist[4][18];
nxt_shortest_dist[4][19] <= shortest_dist[4][19];
nxt_shortest_dist[5][0] <= shortest_dist[5][0];
nxt_shortest_dist[5][1] <= shortest_dist[5][1];
nxt_shortest_dist[5][2] <= shortest_dist[5][2];
nxt_shortest_dist[5][3] <= shortest_dist[5][3];
nxt_shortest_dist[5][4] <= shortest_dist[5][4];
nxt_shortest_dist[5][5] <= shortest_dist[5][5];
nxt_shortest_dist[5][6] <= shortest_dist[5][6];
nxt_shortest_dist[5][7] <= shortest_dist[5][7];
nxt_shortest_dist[5][8] <= shortest_dist[5][8];
nxt_shortest_dist[5][9] <= shortest_dist[5][9];
nxt_shortest_dist[5][10] <= shortest_dist[5][10];
nxt_shortest_dist[5][11] <= shortest_dist[5][11];
nxt_shortest_dist[5][12] <= shortest_dist[5][12];
nxt_shortest_dist[5][13] <= shortest_dist[5][13];
nxt_shortest_dist[5][14] <= shortest_dist[5][14];
nxt_shortest_dist[5][15] <= shortest_dist[5][15];
nxt_shortest_dist[5][16] <= shortest_dist[5][16];
nxt_shortest_dist[5][17] <= shortest_dist[5][17];
nxt_shortest_dist[5][18] <= shortest_dist[5][18];
nxt_shortest_dist[5][19] <= shortest_dist[5][19];
nxt_shortest_dist[6][0] <= shortest_dist[6][0];
nxt_shortest_dist[6][1] <= shortest_dist[6][1];
nxt_shortest_dist[6][2] <= shortest_dist[6][2];
nxt_shortest_dist[6][3] <= shortest_dist[6][3];
nxt_shortest_dist[6][4] <= shortest_dist[6][4];
nxt_shortest_dist[6][5] <= shortest_dist[6][5];
nxt_shortest_dist[6][6] <= shortest_dist[6][6];
nxt_shortest_dist[6][7] <= shortest_dist[6][7];
nxt_shortest_dist[6][8] <= shortest_dist[6][8];
nxt_shortest_dist[6][9] <= shortest_dist[6][9];
nxt_shortest_dist[6][10] <= shortest_dist[6][10];
nxt_shortest_dist[6][11] <= shortest_dist[6][11];
nxt_shortest_dist[6][12] <= shortest_dist[6][12];
nxt_shortest_dist[6][13] <= shortest_dist[6][13];
nxt_shortest_dist[6][14] <= shortest_dist[6][14];
nxt_shortest_dist[6][15] <= shortest_dist[6][15];
nxt_shortest_dist[6][16] <= shortest_dist[6][16];
nxt_shortest_dist[6][17] <= shortest_dist[6][17];
nxt_shortest_dist[6][18] <= shortest_dist[6][18];
nxt_shortest_dist[6][19] <= shortest_dist[6][19];
nxt_shortest_dist[7][0] <= shortest_dist[7][0];
nxt_shortest_dist[7][1] <= shortest_dist[7][1];
nxt_shortest_dist[7][2] <= shortest_dist[7][2];
nxt_shortest_dist[7][3] <= shortest_dist[7][3];
nxt_shortest_dist[7][4] <= shortest_dist[7][4];
nxt_shortest_dist[7][5] <= shortest_dist[7][5];
nxt_shortest_dist[7][6] <= shortest_dist[7][6];
nxt_shortest_dist[7][7] <= shortest_dist[7][7];
nxt_shortest_dist[7][8] <= shortest_dist[7][8];
nxt_shortest_dist[7][9] <= shortest_dist[7][9];
nxt_shortest_dist[7][10] <= shortest_dist[7][10];
nxt_shortest_dist[7][11] <= shortest_dist[7][11];
nxt_shortest_dist[7][12] <= shortest_dist[7][12];
nxt_shortest_dist[7][13] <= shortest_dist[7][13];
nxt_shortest_dist[7][14] <= shortest_dist[7][14];
nxt_shortest_dist[7][15] <= shortest_dist[7][15];
nxt_shortest_dist[7][16] <= shortest_dist[7][16];
nxt_shortest_dist[7][17] <= shortest_dist[7][17];
nxt_shortest_dist[7][18] <= shortest_dist[7][18];
nxt_shortest_dist[7][19] <= shortest_dist[7][19];
nxt_shortest_dist[8][0] <= shortest_dist[8][0];
nxt_shortest_dist[8][1] <= shortest_dist[8][1];
nxt_shortest_dist[8][2] <= shortest_dist[8][2];
nxt_shortest_dist[8][3] <= shortest_dist[8][3];
nxt_shortest_dist[8][4] <= shortest_dist[8][4];
nxt_shortest_dist[8][5] <= shortest_dist[8][5];
nxt_shortest_dist[8][6] <= shortest_dist[8][6];
nxt_shortest_dist[8][7] <= shortest_dist[8][7];
nxt_shortest_dist[8][8] <= shortest_dist[8][8];
nxt_shortest_dist[8][9] <= shortest_dist[8][9];
nxt_shortest_dist[8][10] <= shortest_dist[8][10];
nxt_shortest_dist[8][11] <= shortest_dist[8][11];
nxt_shortest_dist[8][12] <= shortest_dist[8][12];
nxt_shortest_dist[8][13] <= shortest_dist[8][13];
nxt_shortest_dist[8][14] <= shortest_dist[8][14];
nxt_shortest_dist[8][15] <= shortest_dist[8][15];
nxt_shortest_dist[8][16] <= shortest_dist[8][16];
nxt_shortest_dist[8][17] <= shortest_dist[8][17];
nxt_shortest_dist[8][18] <= shortest_dist[8][18];
nxt_shortest_dist[8][19] <= shortest_dist[8][19];
nxt_shortest_dist[9][0] <= shortest_dist[9][0];
nxt_shortest_dist[9][1] <= shortest_dist[9][1];
nxt_shortest_dist[9][2] <= shortest_dist[9][2];
nxt_shortest_dist[9][3] <= shortest_dist[9][3];
nxt_shortest_dist[9][4] <= shortest_dist[9][4];
nxt_shortest_dist[9][5] <= shortest_dist[9][5];
nxt_shortest_dist[9][6] <= shortest_dist[9][6];
nxt_shortest_dist[9][7] <= shortest_dist[9][7];
nxt_shortest_dist[9][8] <= shortest_dist[9][8];
nxt_shortest_dist[9][9] <= shortest_dist[9][9];
nxt_shortest_dist[9][10] <= shortest_dist[9][10];
nxt_shortest_dist[9][11] <= shortest_dist[9][11];
nxt_shortest_dist[9][12] <= shortest_dist[9][12];
nxt_shortest_dist[9][13] <= shortest_dist[9][13];
nxt_shortest_dist[9][14] <= shortest_dist[9][14];
nxt_shortest_dist[9][15] <= shortest_dist[9][15];
nxt_shortest_dist[9][16] <= shortest_dist[9][16];
nxt_shortest_dist[9][17] <= shortest_dist[9][17];
nxt_shortest_dist[9][18] <= shortest_dist[9][18];
nxt_shortest_dist[9][19] <= shortest_dist[9][19];
end
endtask
task bf_init_shortest_path;
begin
nxt_shortest_dist[0][0] <= 1023;
nxt_shortest_dist[0][1] <= 1023;
nxt_shortest_dist[0][2] <= 1023;
nxt_shortest_dist[0][3] <= 1023;
nxt_shortest_dist[0][4] <= 1023;
nxt_shortest_dist[0][5] <= 1023;
nxt_shortest_dist[0][6] <= 1023;
nxt_shortest_dist[0][7] <= 1023;
nxt_shortest_dist[0][8] <= 1023;
nxt_shortest_dist[0][9] <= 1023;
nxt_shortest_dist[0][10] <= 1023;
nxt_shortest_dist[0][11] <= 1023;
nxt_shortest_dist[0][12] <= 1023;
nxt_shortest_dist[0][13] <= 1023;
nxt_shortest_dist[0][14] <= 1023;
nxt_shortest_dist[0][15] <= 1023;
nxt_shortest_dist[0][16] <= 1023;
nxt_shortest_dist[0][17] <= 1023;
nxt_shortest_dist[0][18] <= 1023;
nxt_shortest_dist[0][19] <= 1023;
nxt_shortest_dist[1][0] <= 1023;
nxt_shortest_dist[1][1] <= 1023;
nxt_shortest_dist[1][2] <= 1023;
nxt_shortest_dist[1][3] <= 1023;
nxt_shortest_dist[1][4] <= 1023;
nxt_shortest_dist[1][5] <= 1023;
nxt_shortest_dist[1][6] <= 1023;
nxt_shortest_dist[1][7] <= 1023;
nxt_shortest_dist[1][8] <= 1023;
nxt_shortest_dist[1][9] <= 1023;
nxt_shortest_dist[1][10] <= 1023;
nxt_shortest_dist[1][11] <= 1023;
nxt_shortest_dist[1][12] <= 1023;
nxt_shortest_dist[1][13] <= 1023;
nxt_shortest_dist[1][14] <= 1023;
nxt_shortest_dist[1][15] <= 1023;
nxt_shortest_dist[1][16] <= 1023;
nxt_shortest_dist[1][17] <= 1023;
nxt_shortest_dist[1][18] <= 1023;
nxt_shortest_dist[1][19] <= 1023;
nxt_shortest_dist[2][0] <= 1023;
nxt_shortest_dist[2][1] <= 1023;
nxt_shortest_dist[2][2] <= 1023;
nxt_shortest_dist[2][3] <= 1023;
nxt_shortest_dist[2][4] <= 1023;
nxt_shortest_dist[2][5] <= 1023;
nxt_shortest_dist[2][6] <= 1023;
nxt_shortest_dist[2][7] <= 1023;
nxt_shortest_dist[2][8] <= 1023;
nxt_shortest_dist[2][9] <= 1023;
nxt_shortest_dist[2][10] <= 1023;
nxt_shortest_dist[2][11] <= 1023;
nxt_shortest_dist[2][12] <= 1023;
nxt_shortest_dist[2][13] <= 1023;
nxt_shortest_dist[2][14] <= 1023;
nxt_shortest_dist[2][15] <= 1023;
nxt_shortest_dist[2][16] <= 1023;
nxt_shortest_dist[2][17] <= 1023;
nxt_shortest_dist[2][18] <= 1023;
nxt_shortest_dist[2][19] <= 1023;
nxt_shortest_dist[3][0] <= 1023;
nxt_shortest_dist[3][1] <= 1023;
nxt_shortest_dist[3][2] <= 1023;
nxt_shortest_dist[3][3] <= 1023;
nxt_shortest_dist[3][4] <= 1023;
nxt_shortest_dist[3][5] <= 1023;
nxt_shortest_dist[3][6] <= 1023;
nxt_shortest_dist[3][7] <= 1023;
nxt_shortest_dist[3][8] <= 1023;
nxt_shortest_dist[3][9] <= 1023;
nxt_shortest_dist[3][10] <= 1023;
nxt_shortest_dist[3][11] <= 1023;
nxt_shortest_dist[3][12] <= 1023;
nxt_shortest_dist[3][13] <= 1023;
nxt_shortest_dist[3][14] <= 1023;
nxt_shortest_dist[3][15] <= 1023;
nxt_shortest_dist[3][16] <= 1023;
nxt_shortest_dist[3][17] <= 1023;
nxt_shortest_dist[3][18] <= 1023;
nxt_shortest_dist[3][19] <= 1023;
nxt_shortest_dist[4][0] <= 1023;
nxt_shortest_dist[4][1] <= 1023;
nxt_shortest_dist[4][2] <= 1023;
nxt_shortest_dist[4][3] <= 1023;
nxt_shortest_dist[4][4] <= 1023;
nxt_shortest_dist[4][5] <= 1023;
nxt_shortest_dist[4][6] <= 1023;
nxt_shortest_dist[4][7] <= 1023;
nxt_shortest_dist[4][8] <= 1023;
nxt_shortest_dist[4][9] <= 1023;
nxt_shortest_dist[4][10] <= 1023;
nxt_shortest_dist[4][11] <= 1023;
nxt_shortest_dist[4][12] <= 1023;
nxt_shortest_dist[4][13] <= 1023;
nxt_shortest_dist[4][14] <= 1023;
nxt_shortest_dist[4][15] <= 1023;
nxt_shortest_dist[4][16] <= 1023;
nxt_shortest_dist[4][17] <= 1023;
nxt_shortest_dist[4][18] <= 1023;
nxt_shortest_dist[4][19] <= 1023;
nxt_shortest_dist[5][0] <= 1023;
nxt_shortest_dist[5][1] <= 1023;
nxt_shortest_dist[5][2] <= 1023;
nxt_shortest_dist[5][3] <= 1023;
nxt_shortest_dist[5][4] <= 1023;
nxt_shortest_dist[5][5] <= 1023;
nxt_shortest_dist[5][6] <= 1023;
nxt_shortest_dist[5][7] <= 1023;
nxt_shortest_dist[5][8] <= 1023;
nxt_shortest_dist[5][9] <= 1023;
nxt_shortest_dist[5][10] <= 1023;
nxt_shortest_dist[5][11] <= 1023;
nxt_shortest_dist[5][12] <= 1023;
nxt_shortest_dist[5][13] <= 1023;
nxt_shortest_dist[5][14] <= 1023;
nxt_shortest_dist[5][15] <= 1023;
nxt_shortest_dist[5][16] <= 1023;
nxt_shortest_dist[5][17] <= 1023;
nxt_shortest_dist[5][18] <= 1023;
nxt_shortest_dist[5][19] <= 1023;
nxt_shortest_dist[6][0] <= 1023;
nxt_shortest_dist[6][1] <= 1023;
nxt_shortest_dist[6][2] <= 1023;
nxt_shortest_dist[6][3] <= 1023;
nxt_shortest_dist[6][4] <= 1023;
nxt_shortest_dist[6][5] <= 1023;
nxt_shortest_dist[6][6] <= 1023;
nxt_shortest_dist[6][7] <= 1023;
nxt_shortest_dist[6][8] <= 1023;
nxt_shortest_dist[6][9] <= 1023;
nxt_shortest_dist[6][10] <= 1023;
nxt_shortest_dist[6][11] <= 1023;
nxt_shortest_dist[6][12] <= 1023;
nxt_shortest_dist[6][13] <= 1023;
nxt_shortest_dist[6][14] <= 1023;
nxt_shortest_dist[6][15] <= 1023;
nxt_shortest_dist[6][16] <= 1023;
nxt_shortest_dist[6][17] <= 1023;
nxt_shortest_dist[6][18] <= 1023;
nxt_shortest_dist[6][19] <= 1023;
nxt_shortest_dist[7][0] <= 1023;
nxt_shortest_dist[7][1] <= 1023;
nxt_shortest_dist[7][2] <= 1023;
nxt_shortest_dist[7][3] <= 1023;
nxt_shortest_dist[7][4] <= 1023;
nxt_shortest_dist[7][5] <= 1023;
nxt_shortest_dist[7][6] <= 1023;
nxt_shortest_dist[7][7] <= 1023;
nxt_shortest_dist[7][8] <= 1023;
nxt_shortest_dist[7][9] <= 1023;
nxt_shortest_dist[7][10] <= 1023;
nxt_shortest_dist[7][11] <= 1023;
nxt_shortest_dist[7][12] <= 1023;
nxt_shortest_dist[7][13] <= 1023;
nxt_shortest_dist[7][14] <= 1023;
nxt_shortest_dist[7][15] <= 1023;
nxt_shortest_dist[7][16] <= 1023;
nxt_shortest_dist[7][17] <= 1023;
nxt_shortest_dist[7][18] <= 1023;
nxt_shortest_dist[7][19] <= 1023;
nxt_shortest_dist[8][0] <= 1023;
nxt_shortest_dist[8][1] <= 1023;
nxt_shortest_dist[8][2] <= 1023;
nxt_shortest_dist[8][3] <= 1023;
nxt_shortest_dist[8][4] <= 1023;
nxt_shortest_dist[8][5] <= 1023;
nxt_shortest_dist[8][6] <= 1023;
nxt_shortest_dist[8][7] <= 1023;
nxt_shortest_dist[8][8] <= 1023;
nxt_shortest_dist[8][9] <= 1023;
nxt_shortest_dist[8][10] <= 1023;
nxt_shortest_dist[8][11] <= 1023;
nxt_shortest_dist[8][12] <= 1023;
nxt_shortest_dist[8][13] <= 1023;
nxt_shortest_dist[8][14] <= 1023;
nxt_shortest_dist[8][15] <= 1023;
nxt_shortest_dist[8][16] <= 1023;
nxt_shortest_dist[8][17] <= 1023;
nxt_shortest_dist[8][18] <= 1023;
nxt_shortest_dist[8][19] <= 1023;
nxt_shortest_dist[9][0] <= 1023;
nxt_shortest_dist[9][1] <= 1023;
nxt_shortest_dist[9][2] <= 1023;
nxt_shortest_dist[9][3] <= 1023;
nxt_shortest_dist[9][4] <= 1023;
nxt_shortest_dist[9][5] <= 1023;
nxt_shortest_dist[9][6] <= 1023;
nxt_shortest_dist[9][7] <= 1023;
nxt_shortest_dist[9][8] <= 1023;
nxt_shortest_dist[9][9] <= 1023;
nxt_shortest_dist[9][10] <= 1023;
nxt_shortest_dist[9][11] <= 1023;
nxt_shortest_dist[9][12] <= 1023;
nxt_shortest_dist[9][13] <= 1023;
nxt_shortest_dist[9][14] <= 1023;
nxt_shortest_dist[9][15] <= 1023;
nxt_shortest_dist[9][16] <= 1023;
nxt_shortest_dist[9][17] <= 1023;
nxt_shortest_dist[9][18] <= 1023;
nxt_shortest_dist[9][19] <= 1023;
nxt_shortest_dist[player_r][player_c] <= 0;
end
endtask


	// relax function
	function [2:0] relax_dir;
		input [9:0] ur, uc, dr, dc, lr, lc, rr, rc, original_dist;
		input [2:0] original_dir;
		reg [9:0] tmp, tmp_u, tmp_d, tmp_l, tmp_r;
		reg [2:0] dir, dir_u, dir_d, dir_l, dir_r;
		begin
			tmp = original_dist;
			dir = original_dir;
			tmp_u = (shortest_dist[ur][uc] < tmp-1)? shortest_dist[ur][uc]+1 : tmp;
			dir_u = (shortest_dist[ur][uc] == tmp_u-1)? `MOVE_UP : dir;
			tmp_d = (shortest_dist[dr][dc] < tmp_u-1)? shortest_dist[dr][dc]+1 : tmp_u;
			dir_d = (shortest_dist[dr][dc] == tmp_d-1)? `MOVE_DOWN : dir_u;
			tmp_l = (shortest_dist[lr][lc] < tmp_d-1)? shortest_dist[lr][lc]+1 : tmp_d;
			dir_l = (shortest_dist[lr][lc] == tmp_l-1)? `MOVE_LEFT : dir_d;
			tmp_r = (shortest_dist[rr][rc] < tmp_l-1)? shortest_dist[rr][rc]+1 : tmp_l;
			dir_r = (shortest_dist[rr][rc] == tmp_r-1)? `MOVE_RIGHT : dir_l;
			relax_dir = (tmp_r == 1023)? `MOVE_STOP : dir_r;
		end
	endfunction
	
	function [9:0] relax_dist;
		input [9:0] ur, uc, dr, dc, lr, lc, rr, rc, original_dist;
		reg [9:0] tmp, tmp_u, tmp_d, tmp_l, tmp_r;
		begin
			tmp = original_dist;
			tmp_u = (shortest_dist[ur][uc] < tmp-1)? shortest_dist[ur][uc]+1 : tmp;
			tmp_d = (shortest_dist[dr][dc] < tmp_u-1)? shortest_dist[dr][dc]+1 : tmp_u;
			tmp_l = (shortest_dist[lr][lc] < tmp_d-1)? shortest_dist[lr][lc]+1 : tmp_d;
			tmp_r = (shortest_dist[rr][rc] < tmp_l-1)? shortest_dist[rr][rc]+1 : tmp_l;
			relax_dist = tmp_r;
		end
	endfunction

endmodule